// SPDX-License-Identifier: BSD-2-Clause-Views
/*
 * Copyright (c) 2023 The Regents of the University of California
 */

// Language: Verilog 2001

`resetall
`timescale 1ns / 1ps
`default_nettype none

/*
 * HBM wrapper
 */
module fpga_hbm #
(
    parameter HBM_CH = 32,
    parameter HBM_GROUP_SIZE = HBM_CH,
    parameter AXI_HBM_DATA_WIDTH = 256,
    parameter AXI_HBM_ADDR_WIDTH = 33,
    parameter AXI_HBM_STRB_WIDTH = (AXI_HBM_DATA_WIDTH/8),
    parameter AXI_HBM_ID_WIDTH = 6,
    parameter AXI_HBM_MAX_BURST_LEN = 16
)
(
    input  wire                                  hbm_ref_clk,
    input  wire                                  hbm_rst_in,

    output wire                                  hbm_cattrip_1,
    output wire                                  hbm_cattrip_2,
    output wire [6:0]                            hbm_temp_1,
    output wire [6:0]                            hbm_temp_2,

    output wire [HBM_CH-1:0]                     hbm_clk,
    output wire [HBM_CH-1:0]                     hbm_rst,

    input  wire [HBM_CH*AXI_HBM_ID_WIDTH-1:0]    s_axi_hbm_awid,
    input  wire [HBM_CH*AXI_HBM_ADDR_WIDTH-1:0]  s_axi_hbm_awaddr,
    input  wire [HBM_CH*8-1:0]                   s_axi_hbm_awlen,
    input  wire [HBM_CH*3-1:0]                   s_axi_hbm_awsize,
    input  wire [HBM_CH*2-1:0]                   s_axi_hbm_awburst,
    input  wire [HBM_CH-1:0]                     s_axi_hbm_awlock,
    input  wire [HBM_CH*4-1:0]                   s_axi_hbm_awcache,
    input  wire [HBM_CH*3-1:0]                   s_axi_hbm_awprot,
    input  wire [HBM_CH*4-1:0]                   s_axi_hbm_awqos,
    input  wire [HBM_CH-1:0]                     s_axi_hbm_awvalid,
    output wire [HBM_CH-1:0]                     s_axi_hbm_awready,
    input  wire [HBM_CH*AXI_HBM_DATA_WIDTH-1:0]  s_axi_hbm_wdata,
    input  wire [HBM_CH*AXI_HBM_STRB_WIDTH-1:0]  s_axi_hbm_wstrb,
    input  wire [HBM_CH-1:0]                     s_axi_hbm_wlast,
    input  wire [HBM_CH-1:0]                     s_axi_hbm_wvalid,
    output wire [HBM_CH-1:0]                     s_axi_hbm_wready,
    output wire [HBM_CH*AXI_HBM_ID_WIDTH-1:0]    s_axi_hbm_bid,
    output wire [HBM_CH*2-1:0]                   s_axi_hbm_bresp,
    output wire [HBM_CH-1:0]                     s_axi_hbm_bvalid,
    input  wire [HBM_CH-1:0]                     s_axi_hbm_bready,
    input  wire [HBM_CH*AXI_HBM_ID_WIDTH-1:0]    s_axi_hbm_arid,
    input  wire [HBM_CH*AXI_HBM_ADDR_WIDTH-1:0]  s_axi_hbm_araddr,
    input  wire [HBM_CH*8-1:0]                   s_axi_hbm_arlen,
    input  wire [HBM_CH*3-1:0]                   s_axi_hbm_arsize,
    input  wire [HBM_CH*2-1:0]                   s_axi_hbm_arburst,
    input  wire [HBM_CH-1:0]                     s_axi_hbm_arlock,
    input  wire [HBM_CH*4-1:0]                   s_axi_hbm_arcache,
    input  wire [HBM_CH*3-1:0]                   s_axi_hbm_arprot,
    input  wire [HBM_CH*4-1:0]                   s_axi_hbm_arqos,
    input  wire [HBM_CH-1:0]                     s_axi_hbm_arvalid,
    output wire [HBM_CH-1:0]                     s_axi_hbm_arready,
    output wire [HBM_CH*AXI_HBM_ID_WIDTH-1:0]    s_axi_hbm_rid,
    output wire [HBM_CH*AXI_HBM_DATA_WIDTH-1:0]  s_axi_hbm_rdata,
    output wire [HBM_CH*2-1:0]                   s_axi_hbm_rresp,
    output wire [HBM_CH-1:0]                     s_axi_hbm_rlast,
    output wire [HBM_CH-1:0]                     s_axi_hbm_rvalid,
    input  wire [HBM_CH-1:0]                     s_axi_hbm_rready,

    output wire [HBM_CH-1:0]                     hbm_status
);

localparam HBM_CH_INT = 32;
localparam HBM_CH_STRIDE = HBM_CH_INT / 2**$clog2(HBM_CH);

wire [HBM_CH_INT-1:0]                     hbm_clk_int;
wire [HBM_CH_INT-1:0]                     hbm_rst_int;

wire [HBM_CH_INT*AXI_HBM_ID_WIDTH-1:0]    m_axi_hbm_int_awid;
wire [HBM_CH_INT*AXI_HBM_ADDR_WIDTH-1:0]  m_axi_hbm_int_awaddr;
wire [HBM_CH_INT*8-1:0]                   m_axi_hbm_int_awlen;
wire [HBM_CH_INT*3-1:0]                   m_axi_hbm_int_awsize;
wire [HBM_CH_INT*2-1:0]                   m_axi_hbm_int_awburst;
wire [HBM_CH_INT-1:0]                     m_axi_hbm_int_awlock;
wire [HBM_CH_INT*4-1:0]                   m_axi_hbm_int_awcache;
wire [HBM_CH_INT*3-1:0]                   m_axi_hbm_int_awprot;
wire [HBM_CH_INT*4-1:0]                   m_axi_hbm_int_awqos;
wire [HBM_CH_INT-1:0]                     m_axi_hbm_int_awvalid;
wire [HBM_CH_INT-1:0]                     m_axi_hbm_int_awready;
wire [HBM_CH_INT*AXI_HBM_DATA_WIDTH-1:0]  m_axi_hbm_int_wdata;
wire [HBM_CH_INT*AXI_HBM_STRB_WIDTH-1:0]  m_axi_hbm_int_wstrb;
wire [HBM_CH_INT-1:0]                     m_axi_hbm_int_wlast;
wire [HBM_CH_INT-1:0]                     m_axi_hbm_int_wvalid;
wire [HBM_CH_INT-1:0]                     m_axi_hbm_int_wready;
wire [HBM_CH_INT*AXI_HBM_ID_WIDTH-1:0]    m_axi_hbm_int_bid;
wire [HBM_CH_INT*2-1:0]                   m_axi_hbm_int_bresp;
wire [HBM_CH_INT-1:0]                     m_axi_hbm_int_bvalid;
wire [HBM_CH_INT-1:0]                     m_axi_hbm_int_bready;
wire [HBM_CH_INT*AXI_HBM_ID_WIDTH-1:0]    m_axi_hbm_int_arid;
wire [HBM_CH_INT*AXI_HBM_ADDR_WIDTH-1:0]  m_axi_hbm_int_araddr;
wire [HBM_CH_INT*8-1:0]                   m_axi_hbm_int_arlen;
wire [HBM_CH_INT*3-1:0]                   m_axi_hbm_int_arsize;
wire [HBM_CH_INT*2-1:0]                   m_axi_hbm_int_arburst;
wire [HBM_CH_INT-1:0]                     m_axi_hbm_int_arlock;
wire [HBM_CH_INT*4-1:0]                   m_axi_hbm_int_arcache;
wire [HBM_CH_INT*3-1:0]                   m_axi_hbm_int_arprot;
wire [HBM_CH_INT*4-1:0]                   m_axi_hbm_int_arqos;
wire [HBM_CH_INT-1:0]                     m_axi_hbm_int_arvalid;
wire [HBM_CH_INT-1:0]                     m_axi_hbm_int_arready;
wire [HBM_CH_INT*AXI_HBM_ID_WIDTH-1:0]    m_axi_hbm_int_rid;
wire [HBM_CH_INT*AXI_HBM_DATA_WIDTH-1:0]  m_axi_hbm_int_rdata;
wire [HBM_CH_INT*2-1:0]                   m_axi_hbm_int_rresp;
wire [HBM_CH_INT-1:0]                     m_axi_hbm_int_rlast;
wire [HBM_CH_INT-1:0]                     m_axi_hbm_int_rvalid;
wire [HBM_CH_INT-1:0]                     m_axi_hbm_int_rready;

generate

genvar n;

wire hbm_mmcm_rst = hbm_rst_in;
wire hbm_mmcm_locked;
wire hbm_mmcm_clkfb;

wire hbm_axi_clk_mmcm;
wire hbm_axi_clk;
wire hbm_axi_rst_int;
wire hbm_axi_rst;

// HBM MMCM instance
// 100 MHz in, 450 MHz out
// PFD range: 10 MHz to 500 MHz
// VCO range: 800 MHz to 1600 MHz
// M = 9, D = 1 sets Fvco = 900 MHz
// Divide by 2 to get output frequency of 450 MHz
MMCME4_BASE #(
    .BANDWIDTH("OPTIMIZED"),
    .CLKOUT0_DIVIDE_F(2),
    .CLKOUT0_DUTY_CYCLE(0.5),
    .CLKOUT0_PHASE(0),
    .CLKOUT1_DIVIDE(1),
    .CLKOUT1_DUTY_CYCLE(0.5),
    .CLKOUT1_PHASE(0),
    .CLKOUT2_DIVIDE(1),
    .CLKOUT2_DUTY_CYCLE(0.5),
    .CLKOUT2_PHASE(0),
    .CLKOUT3_DIVIDE(1),
    .CLKOUT3_DUTY_CYCLE(0.5),
    .CLKOUT3_PHASE(0),
    .CLKOUT4_DIVIDE(1),
    .CLKOUT4_DUTY_CYCLE(0.5),
    .CLKOUT4_PHASE(0),
    .CLKOUT5_DIVIDE(1),
    .CLKOUT5_DUTY_CYCLE(0.5),
    .CLKOUT5_PHASE(0),
    .CLKOUT6_DIVIDE(1),
    .CLKOUT6_DUTY_CYCLE(0.5),
    .CLKOUT6_PHASE(0),
    .CLKFBOUT_MULT_F(9),
    .CLKFBOUT_PHASE(0),
    .DIVCLK_DIVIDE(1),
    .REF_JITTER1(0.010),
    .CLKIN1_PERIOD(10.000),
    .STARTUP_WAIT("FALSE"),
    .CLKOUT4_CASCADE("FALSE")
)
hbm_mmcm_inst (
    .CLKIN1(hbm_ref_clk),
    .CLKFBIN(hbm_mmcm_clkfb),
    .RST(hbm_mmcm_rst),
    .PWRDWN(1'b0),
    .CLKOUT0(hbm_axi_clk_mmcm),
    .CLKOUT0B(),
    .CLKOUT1(),
    .CLKOUT1B(),
    .CLKOUT2(),
    .CLKOUT2B(),
    .CLKOUT3(),
    .CLKOUT3B(),
    .CLKOUT4(),
    .CLKOUT5(),
    .CLKOUT6(),
    .CLKFBOUT(hbm_mmcm_clkfb),
    .CLKFBOUTB(),
    .LOCKED(hbm_mmcm_locked)
);

BUFG
hbm_axi_clk_bufg_inst (
    .I(hbm_axi_clk_mmcm),
    .O(hbm_axi_clk)
);

sync_reset #(
    .N(4)
)
sync_reset_hbm_axi_inst (
    .clk(hbm_axi_clk),
    .rst(~hbm_mmcm_locked),
    .out(hbm_axi_rst_int)
);

// extra register for hbm_axi_rst signal
(* shreg_extract = "no" *)
reg hbm_axi_rst_reg_1 = 1'b1;
(* shreg_extract = "no" *)
reg hbm_axi_rst_reg_2 = 1'b1;

always @(posedge hbm_axi_clk) begin
    hbm_axi_rst_reg_1 <= hbm_axi_rst_int;
    hbm_axi_rst_reg_2 <= hbm_axi_rst_reg_1;
end

BUFG
hbm_axi_rst_bufg_inst (
    .I(hbm_axi_rst_reg_2),
    .O(hbm_axi_rst)
);

assign hbm_clk_int = {HBM_CH_INT{hbm_axi_clk}};
assign hbm_rst_int = {HBM_CH_INT{hbm_axi_rst}};

hbm_0 hbm_inst (
    .HBM_REF_CLK_0(hbm_ref_clk),
    .HBM_REF_CLK_1(hbm_ref_clk),

    .APB_0_PWDATA(32'd0),
    .APB_0_PADDR(22'd0),
    .APB_0_PCLK(hbm_ref_clk),
    .APB_0_PENABLE(1'b0),
    .APB_0_PRESET_N(1'b1),
    .APB_0_PSEL(1'b0),
    .APB_0_PWRITE(1'b0),
    .APB_0_PRDATA(),
    .APB_0_PREADY(),
    .APB_0_PSLVERR(),
    .apb_complete_0(),

    .APB_1_PWDATA(32'd0),
    .APB_1_PADDR(22'd0),
    .APB_1_PCLK(hbm_ref_clk),
    .APB_1_PENABLE(1'b0),
    .APB_1_PRESET_N(1'b1),
    .APB_1_PSEL(1'b0),
    .APB_1_PWRITE(1'b0),
    .APB_1_PRDATA(),
    .APB_1_PREADY(),
    .APB_1_PSLVERR(),
    .apb_complete_1(),

    .AXI_00_ACLK(hbm_clk_int[0 +: 1]),
    .AXI_00_ARESET_N(!hbm_rst_int[0 +: 1]),

    .AXI_00_ARADDR(m_axi_hbm_int_araddr[0*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_00_ARBURST(m_axi_hbm_int_arburst[0*2 +: 2]),
    .AXI_00_ARID(m_axi_hbm_int_arid[0*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_00_ARLEN(m_axi_hbm_int_arlen[0*8 +: 4]),
    .AXI_00_ARSIZE(m_axi_hbm_int_arsize[0*3 +: 3]),
    .AXI_00_ARVALID(m_axi_hbm_int_arvalid[0 +: 1]),
    .AXI_00_ARREADY(m_axi_hbm_int_arready[0 +: 1]),
    .AXI_00_RDATA_PARITY(),
    .AXI_00_RDATA(m_axi_hbm_int_rdata[0*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_00_RID(m_axi_hbm_int_rid[0*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_00_RLAST(m_axi_hbm_int_rlast[0 +: 1]),
    .AXI_00_RRESP(m_axi_hbm_int_rresp[0*2 +: 2]),
    .AXI_00_RVALID(m_axi_hbm_int_rvalid[0 +: 1]),
    .AXI_00_RREADY(m_axi_hbm_int_rready[0 +: 1]),
    .AXI_00_AWADDR(m_axi_hbm_int_awaddr[0*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_00_AWBURST(m_axi_hbm_int_awburst[0*2 +: 2]),
    .AXI_00_AWID(m_axi_hbm_int_awid[0*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_00_AWLEN(m_axi_hbm_int_awlen[0*8 +: 4]),
    .AXI_00_AWSIZE(m_axi_hbm_int_awsize[0*3 +: 3]),
    .AXI_00_AWVALID(m_axi_hbm_int_awvalid[0 +: 1]),
    .AXI_00_AWREADY(m_axi_hbm_int_awready[0 +: 1]),
    .AXI_00_WDATA(m_axi_hbm_int_wdata[0*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_00_WLAST(m_axi_hbm_int_wlast[0 +: 1]),
    .AXI_00_WSTRB(m_axi_hbm_int_wstrb[0*AXI_HBM_STRB_WIDTH +: AXI_HBM_STRB_WIDTH]),
    .AXI_00_WDATA_PARITY(32'd0),
    .AXI_00_WVALID(m_axi_hbm_int_wvalid[0 +: 1]),
    .AXI_00_WREADY(m_axi_hbm_int_wready[0 +: 1]),
    .AXI_00_BID(m_axi_hbm_int_bid[0*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_00_BRESP(m_axi_hbm_int_bresp[0*2 +: 2]),
    .AXI_00_BVALID(m_axi_hbm_int_bvalid[0 +: 1]),
    .AXI_00_BREADY(m_axi_hbm_int_bready[0 +: 1]),

    .AXI_01_ACLK(hbm_clk_int[1 +: 1]),
    .AXI_01_ARESET_N(!hbm_rst_int[1 +: 1]),

    .AXI_01_ARADDR(m_axi_hbm_int_araddr[1*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_01_ARBURST(m_axi_hbm_int_arburst[1*2 +: 2]),
    .AXI_01_ARID(m_axi_hbm_int_arid[1*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_01_ARLEN(m_axi_hbm_int_arlen[1*8 +: 4]),
    .AXI_01_ARSIZE(m_axi_hbm_int_arsize[1*3 +: 3]),
    .AXI_01_ARVALID(m_axi_hbm_int_arvalid[1 +: 1]),
    .AXI_01_ARREADY(m_axi_hbm_int_arready[1 +: 1]),
    .AXI_01_RDATA_PARITY(),
    .AXI_01_RDATA(m_axi_hbm_int_rdata[1*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_01_RID(m_axi_hbm_int_rid[1*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_01_RLAST(m_axi_hbm_int_rlast[1 +: 1]),
    .AXI_01_RRESP(m_axi_hbm_int_rresp[1*2 +: 2]),
    .AXI_01_RVALID(m_axi_hbm_int_rvalid[1 +: 1]),
    .AXI_01_RREADY(m_axi_hbm_int_rready[1 +: 1]),
    .AXI_01_AWADDR(m_axi_hbm_int_awaddr[1*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_01_AWBURST(m_axi_hbm_int_awburst[1*2 +: 2]),
    .AXI_01_AWID(m_axi_hbm_int_awid[1*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_01_AWLEN(m_axi_hbm_int_awlen[1*8 +: 4]),
    .AXI_01_AWSIZE(m_axi_hbm_int_awsize[1*3 +: 3]),
    .AXI_01_AWVALID(m_axi_hbm_int_awvalid[1 +: 1]),
    .AXI_01_AWREADY(m_axi_hbm_int_awready[1 +: 1]),
    .AXI_01_WDATA(m_axi_hbm_int_wdata[1*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_01_WLAST(m_axi_hbm_int_wlast[1 +: 1]),
    .AXI_01_WSTRB(m_axi_hbm_int_wstrb[1*AXI_HBM_STRB_WIDTH +: AXI_HBM_STRB_WIDTH]),
    .AXI_01_WDATA_PARITY(32'd0),
    .AXI_01_WVALID(m_axi_hbm_int_wvalid[1 +: 1]),
    .AXI_01_WREADY(m_axi_hbm_int_wready[1 +: 1]),
    .AXI_01_BID(m_axi_hbm_int_bid[1*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_01_BRESP(m_axi_hbm_int_bresp[1*2 +: 2]),
    .AXI_01_BVALID(m_axi_hbm_int_bvalid[1 +: 1]),
    .AXI_01_BREADY(m_axi_hbm_int_bready[1 +: 1]),

    .AXI_02_ACLK(hbm_clk_int[2 +: 1]),
    .AXI_02_ARESET_N(!hbm_rst_int[2 +: 1]),

    .AXI_02_ARADDR(m_axi_hbm_int_araddr[2*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_02_ARBURST(m_axi_hbm_int_arburst[2*2 +: 2]),
    .AXI_02_ARID(m_axi_hbm_int_arid[2*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_02_ARLEN(m_axi_hbm_int_arlen[2*8 +: 4]),
    .AXI_02_ARSIZE(m_axi_hbm_int_arsize[2*3 +: 3]),
    .AXI_02_ARVALID(m_axi_hbm_int_arvalid[2 +: 1]),
    .AXI_02_ARREADY(m_axi_hbm_int_arready[2 +: 1]),
    .AXI_02_RDATA_PARITY(),
    .AXI_02_RDATA(m_axi_hbm_int_rdata[2*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_02_RID(m_axi_hbm_int_rid[2*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_02_RLAST(m_axi_hbm_int_rlast[2 +: 1]),
    .AXI_02_RRESP(m_axi_hbm_int_rresp[2*2 +: 2]),
    .AXI_02_RVALID(m_axi_hbm_int_rvalid[2 +: 1]),
    .AXI_02_RREADY(m_axi_hbm_int_rready[2 +: 1]),
    .AXI_02_AWADDR(m_axi_hbm_int_awaddr[2*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_02_AWBURST(m_axi_hbm_int_awburst[2*2 +: 2]),
    .AXI_02_AWID(m_axi_hbm_int_awid[2*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_02_AWLEN(m_axi_hbm_int_awlen[2*8 +: 4]),
    .AXI_02_AWSIZE(m_axi_hbm_int_awsize[2*3 +: 3]),
    .AXI_02_AWVALID(m_axi_hbm_int_awvalid[2 +: 1]),
    .AXI_02_AWREADY(m_axi_hbm_int_awready[2 +: 1]),
    .AXI_02_WDATA(m_axi_hbm_int_wdata[2*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_02_WLAST(m_axi_hbm_int_wlast[2 +: 1]),
    .AXI_02_WSTRB(m_axi_hbm_int_wstrb[2*AXI_HBM_STRB_WIDTH +: AXI_HBM_STRB_WIDTH]),
    .AXI_02_WDATA_PARITY(32'd0),
    .AXI_02_WVALID(m_axi_hbm_int_wvalid[2 +: 1]),
    .AXI_02_WREADY(m_axi_hbm_int_wready[2 +: 1]),
    .AXI_02_BID(m_axi_hbm_int_bid[2*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_02_BRESP(m_axi_hbm_int_bresp[2*2 +: 2]),
    .AXI_02_BVALID(m_axi_hbm_int_bvalid[2 +: 1]),
    .AXI_02_BREADY(m_axi_hbm_int_bready[2 +: 1]),

    .AXI_03_ACLK(hbm_clk_int[3 +: 1]),
    .AXI_03_ARESET_N(!hbm_rst_int[3 +: 1]),

    .AXI_03_ARADDR(m_axi_hbm_int_araddr[3*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_03_ARBURST(m_axi_hbm_int_arburst[3*2 +: 2]),
    .AXI_03_ARID(m_axi_hbm_int_arid[3*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_03_ARLEN(m_axi_hbm_int_arlen[3*8 +: 4]),
    .AXI_03_ARSIZE(m_axi_hbm_int_arsize[3*3 +: 3]),
    .AXI_03_ARVALID(m_axi_hbm_int_arvalid[3 +: 1]),
    .AXI_03_ARREADY(m_axi_hbm_int_arready[3 +: 1]),
    .AXI_03_RDATA_PARITY(),
    .AXI_03_RDATA(m_axi_hbm_int_rdata[3*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_03_RID(m_axi_hbm_int_rid[3*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_03_RLAST(m_axi_hbm_int_rlast[3 +: 1]),
    .AXI_03_RRESP(m_axi_hbm_int_rresp[3*2 +: 2]),
    .AXI_03_RVALID(m_axi_hbm_int_rvalid[3 +: 1]),
    .AXI_03_RREADY(m_axi_hbm_int_rready[3 +: 1]),
    .AXI_03_AWADDR(m_axi_hbm_int_awaddr[3*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_03_AWBURST(m_axi_hbm_int_awburst[3*2 +: 2]),
    .AXI_03_AWID(m_axi_hbm_int_awid[3*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_03_AWLEN(m_axi_hbm_int_awlen[3*8 +: 4]),
    .AXI_03_AWSIZE(m_axi_hbm_int_awsize[3*3 +: 3]),
    .AXI_03_AWVALID(m_axi_hbm_int_awvalid[3 +: 1]),
    .AXI_03_AWREADY(m_axi_hbm_int_awready[3 +: 1]),
    .AXI_03_WDATA(m_axi_hbm_int_wdata[3*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_03_WLAST(m_axi_hbm_int_wlast[3 +: 1]),
    .AXI_03_WSTRB(m_axi_hbm_int_wstrb[3*AXI_HBM_STRB_WIDTH +: AXI_HBM_STRB_WIDTH]),
    .AXI_03_WDATA_PARITY(32'd0),
    .AXI_03_WVALID(m_axi_hbm_int_wvalid[3 +: 1]),
    .AXI_03_WREADY(m_axi_hbm_int_wready[3 +: 1]),
    .AXI_03_BID(m_axi_hbm_int_bid[3*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_03_BRESP(m_axi_hbm_int_bresp[3*2 +: 2]),
    .AXI_03_BVALID(m_axi_hbm_int_bvalid[3 +: 1]),
    .AXI_03_BREADY(m_axi_hbm_int_bready[3 +: 1]),

    .AXI_04_ACLK(hbm_clk_int[4 +: 1]),
    .AXI_04_ARESET_N(!hbm_rst_int[4 +: 1]),

    .AXI_04_ARADDR(m_axi_hbm_int_araddr[4*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_04_ARBURST(m_axi_hbm_int_arburst[4*2 +: 2]),
    .AXI_04_ARID(m_axi_hbm_int_arid[4*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_04_ARLEN(m_axi_hbm_int_arlen[4*8 +: 4]),
    .AXI_04_ARSIZE(m_axi_hbm_int_arsize[4*3 +: 3]),
    .AXI_04_ARVALID(m_axi_hbm_int_arvalid[4 +: 1]),
    .AXI_04_ARREADY(m_axi_hbm_int_arready[4 +: 1]),
    .AXI_04_RDATA_PARITY(),
    .AXI_04_RDATA(m_axi_hbm_int_rdata[4*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_04_RID(m_axi_hbm_int_rid[4*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_04_RLAST(m_axi_hbm_int_rlast[4 +: 1]),
    .AXI_04_RRESP(m_axi_hbm_int_rresp[4*2 +: 2]),
    .AXI_04_RVALID(m_axi_hbm_int_rvalid[4 +: 1]),
    .AXI_04_RREADY(m_axi_hbm_int_rready[4 +: 1]),
    .AXI_04_AWADDR(m_axi_hbm_int_awaddr[4*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_04_AWBURST(m_axi_hbm_int_awburst[4*2 +: 2]),
    .AXI_04_AWID(m_axi_hbm_int_awid[4*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_04_AWLEN(m_axi_hbm_int_awlen[4*8 +: 4]),
    .AXI_04_AWSIZE(m_axi_hbm_int_awsize[4*3 +: 3]),
    .AXI_04_AWVALID(m_axi_hbm_int_awvalid[4 +: 1]),
    .AXI_04_AWREADY(m_axi_hbm_int_awready[4 +: 1]),
    .AXI_04_WDATA(m_axi_hbm_int_wdata[4*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_04_WLAST(m_axi_hbm_int_wlast[4 +: 1]),
    .AXI_04_WSTRB(m_axi_hbm_int_wstrb[4*AXI_HBM_STRB_WIDTH +: AXI_HBM_STRB_WIDTH]),
    .AXI_04_WDATA_PARITY(32'd0),
    .AXI_04_WVALID(m_axi_hbm_int_wvalid[4 +: 1]),
    .AXI_04_WREADY(m_axi_hbm_int_wready[4 +: 1]),
    .AXI_04_BID(m_axi_hbm_int_bid[4*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_04_BRESP(m_axi_hbm_int_bresp[4*2 +: 2]),
    .AXI_04_BVALID(m_axi_hbm_int_bvalid[4 +: 1]),
    .AXI_04_BREADY(m_axi_hbm_int_bready[4 +: 1]),

    .AXI_05_ACLK(hbm_clk_int[5 +: 1]),
    .AXI_05_ARESET_N(!hbm_rst_int[5 +: 1]),

    .AXI_05_ARADDR(m_axi_hbm_int_araddr[5*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_05_ARBURST(m_axi_hbm_int_arburst[5*2 +: 2]),
    .AXI_05_ARID(m_axi_hbm_int_arid[5*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_05_ARLEN(m_axi_hbm_int_arlen[5*8 +: 4]),
    .AXI_05_ARSIZE(m_axi_hbm_int_arsize[5*3 +: 3]),
    .AXI_05_ARVALID(m_axi_hbm_int_arvalid[5 +: 1]),
    .AXI_05_ARREADY(m_axi_hbm_int_arready[5 +: 1]),
    .AXI_05_RDATA_PARITY(),
    .AXI_05_RDATA(m_axi_hbm_int_rdata[5*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_05_RID(m_axi_hbm_int_rid[5*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_05_RLAST(m_axi_hbm_int_rlast[5 +: 1]),
    .AXI_05_RRESP(m_axi_hbm_int_rresp[5*2 +: 2]),
    .AXI_05_RVALID(m_axi_hbm_int_rvalid[5 +: 1]),
    .AXI_05_RREADY(m_axi_hbm_int_rready[5 +: 1]),
    .AXI_05_AWADDR(m_axi_hbm_int_awaddr[5*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_05_AWBURST(m_axi_hbm_int_awburst[5*2 +: 2]),
    .AXI_05_AWID(m_axi_hbm_int_awid[5*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_05_AWLEN(m_axi_hbm_int_awlen[5*8 +: 4]),
    .AXI_05_AWSIZE(m_axi_hbm_int_awsize[5*3 +: 3]),
    .AXI_05_AWVALID(m_axi_hbm_int_awvalid[5 +: 1]),
    .AXI_05_AWREADY(m_axi_hbm_int_awready[5 +: 1]),
    .AXI_05_WDATA(m_axi_hbm_int_wdata[5*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_05_WLAST(m_axi_hbm_int_wlast[5 +: 1]),
    .AXI_05_WSTRB(m_axi_hbm_int_wstrb[5*AXI_HBM_STRB_WIDTH +: AXI_HBM_STRB_WIDTH]),
    .AXI_05_WDATA_PARITY(32'd0),
    .AXI_05_WVALID(m_axi_hbm_int_wvalid[5 +: 1]),
    .AXI_05_WREADY(m_axi_hbm_int_wready[5 +: 1]),
    .AXI_05_BID(m_axi_hbm_int_bid[5*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_05_BRESP(m_axi_hbm_int_bresp[5*2 +: 2]),
    .AXI_05_BVALID(m_axi_hbm_int_bvalid[5 +: 1]),
    .AXI_05_BREADY(m_axi_hbm_int_bready[5 +: 1]),

    .AXI_06_ACLK(hbm_clk_int[6 +: 1]),
    .AXI_06_ARESET_N(!hbm_rst_int[6 +: 1]),

    .AXI_06_ARADDR(m_axi_hbm_int_araddr[6*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_06_ARBURST(m_axi_hbm_int_arburst[6*2 +: 2]),
    .AXI_06_ARID(m_axi_hbm_int_arid[6*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_06_ARLEN(m_axi_hbm_int_arlen[6*8 +: 4]),
    .AXI_06_ARSIZE(m_axi_hbm_int_arsize[6*3 +: 3]),
    .AXI_06_ARVALID(m_axi_hbm_int_arvalid[6 +: 1]),
    .AXI_06_ARREADY(m_axi_hbm_int_arready[6 +: 1]),
    .AXI_06_RDATA_PARITY(),
    .AXI_06_RDATA(m_axi_hbm_int_rdata[6*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_06_RID(m_axi_hbm_int_rid[6*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_06_RLAST(m_axi_hbm_int_rlast[6 +: 1]),
    .AXI_06_RRESP(m_axi_hbm_int_rresp[6*2 +: 2]),
    .AXI_06_RVALID(m_axi_hbm_int_rvalid[6 +: 1]),
    .AXI_06_RREADY(m_axi_hbm_int_rready[6 +: 1]),
    .AXI_06_AWADDR(m_axi_hbm_int_awaddr[6*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_06_AWBURST(m_axi_hbm_int_awburst[6*2 +: 2]),
    .AXI_06_AWID(m_axi_hbm_int_awid[6*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_06_AWLEN(m_axi_hbm_int_awlen[6*8 +: 4]),
    .AXI_06_AWSIZE(m_axi_hbm_int_awsize[6*3 +: 3]),
    .AXI_06_AWVALID(m_axi_hbm_int_awvalid[6 +: 1]),
    .AXI_06_AWREADY(m_axi_hbm_int_awready[6 +: 1]),
    .AXI_06_WDATA(m_axi_hbm_int_wdata[6*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_06_WLAST(m_axi_hbm_int_wlast[6 +: 1]),
    .AXI_06_WSTRB(m_axi_hbm_int_wstrb[6*AXI_HBM_STRB_WIDTH +: AXI_HBM_STRB_WIDTH]),
    .AXI_06_WDATA_PARITY(32'd0),
    .AXI_06_WVALID(m_axi_hbm_int_wvalid[6 +: 1]),
    .AXI_06_WREADY(m_axi_hbm_int_wready[6 +: 1]),
    .AXI_06_BID(m_axi_hbm_int_bid[6*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_06_BRESP(m_axi_hbm_int_bresp[6*2 +: 2]),
    .AXI_06_BVALID(m_axi_hbm_int_bvalid[6 +: 1]),
    .AXI_06_BREADY(m_axi_hbm_int_bready[6 +: 1]),

    .AXI_07_ACLK(hbm_clk_int[7 +: 1]),
    .AXI_07_ARESET_N(!hbm_rst_int[7 +: 1]),

    .AXI_07_ARADDR(m_axi_hbm_int_araddr[7*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_07_ARBURST(m_axi_hbm_int_arburst[7*2 +: 2]),
    .AXI_07_ARID(m_axi_hbm_int_arid[7*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_07_ARLEN(m_axi_hbm_int_arlen[7*8 +: 4]),
    .AXI_07_ARSIZE(m_axi_hbm_int_arsize[7*3 +: 3]),
    .AXI_07_ARVALID(m_axi_hbm_int_arvalid[7 +: 1]),
    .AXI_07_ARREADY(m_axi_hbm_int_arready[7 +: 1]),
    .AXI_07_RDATA_PARITY(),
    .AXI_07_RDATA(m_axi_hbm_int_rdata[7*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_07_RID(m_axi_hbm_int_rid[7*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_07_RLAST(m_axi_hbm_int_rlast[7 +: 1]),
    .AXI_07_RRESP(m_axi_hbm_int_rresp[7*2 +: 2]),
    .AXI_07_RVALID(m_axi_hbm_int_rvalid[7 +: 1]),
    .AXI_07_RREADY(m_axi_hbm_int_rready[7 +: 1]),
    .AXI_07_AWADDR(m_axi_hbm_int_awaddr[7*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_07_AWBURST(m_axi_hbm_int_awburst[7*2 +: 2]),
    .AXI_07_AWID(m_axi_hbm_int_awid[7*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_07_AWLEN(m_axi_hbm_int_awlen[7*8 +: 4]),
    .AXI_07_AWSIZE(m_axi_hbm_int_awsize[7*3 +: 3]),
    .AXI_07_AWVALID(m_axi_hbm_int_awvalid[7 +: 1]),
    .AXI_07_AWREADY(m_axi_hbm_int_awready[7 +: 1]),
    .AXI_07_WDATA(m_axi_hbm_int_wdata[7*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_07_WLAST(m_axi_hbm_int_wlast[7 +: 1]),
    .AXI_07_WSTRB(m_axi_hbm_int_wstrb[7*AXI_HBM_STRB_WIDTH +: AXI_HBM_STRB_WIDTH]),
    .AXI_07_WDATA_PARITY(32'd0),
    .AXI_07_WVALID(m_axi_hbm_int_wvalid[7 +: 1]),
    .AXI_07_WREADY(m_axi_hbm_int_wready[7 +: 1]),
    .AXI_07_BID(m_axi_hbm_int_bid[7*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_07_BRESP(m_axi_hbm_int_bresp[7*2 +: 2]),
    .AXI_07_BVALID(m_axi_hbm_int_bvalid[7 +: 1]),
    .AXI_07_BREADY(m_axi_hbm_int_bready[7 +: 1]),

    .AXI_08_ACLK(hbm_clk_int[8 +: 1]),
    .AXI_08_ARESET_N(!hbm_rst_int[8 +: 1]),

    .AXI_08_ARADDR(m_axi_hbm_int_araddr[8*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_08_ARBURST(m_axi_hbm_int_arburst[8*2 +: 2]),
    .AXI_08_ARID(m_axi_hbm_int_arid[8*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_08_ARLEN(m_axi_hbm_int_arlen[8*8 +: 4]),
    .AXI_08_ARSIZE(m_axi_hbm_int_arsize[8*3 +: 3]),
    .AXI_08_ARVALID(m_axi_hbm_int_arvalid[8 +: 1]),
    .AXI_08_ARREADY(m_axi_hbm_int_arready[8 +: 1]),
    .AXI_08_RDATA_PARITY(),
    .AXI_08_RDATA(m_axi_hbm_int_rdata[8*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_08_RID(m_axi_hbm_int_rid[8*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_08_RLAST(m_axi_hbm_int_rlast[8 +: 1]),
    .AXI_08_RRESP(m_axi_hbm_int_rresp[8*2 +: 2]),
    .AXI_08_RVALID(m_axi_hbm_int_rvalid[8 +: 1]),
    .AXI_08_RREADY(m_axi_hbm_int_rready[8 +: 1]),
    .AXI_08_AWADDR(m_axi_hbm_int_awaddr[8*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_08_AWBURST(m_axi_hbm_int_awburst[8*2 +: 2]),
    .AXI_08_AWID(m_axi_hbm_int_awid[8*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_08_AWLEN(m_axi_hbm_int_awlen[8*8 +: 4]),
    .AXI_08_AWSIZE(m_axi_hbm_int_awsize[8*3 +: 3]),
    .AXI_08_AWVALID(m_axi_hbm_int_awvalid[8 +: 1]),
    .AXI_08_AWREADY(m_axi_hbm_int_awready[8 +: 1]),
    .AXI_08_WDATA(m_axi_hbm_int_wdata[8*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_08_WLAST(m_axi_hbm_int_wlast[8 +: 1]),
    .AXI_08_WSTRB(m_axi_hbm_int_wstrb[8*AXI_HBM_STRB_WIDTH +: AXI_HBM_STRB_WIDTH]),
    .AXI_08_WDATA_PARITY(32'd0),
    .AXI_08_WVALID(m_axi_hbm_int_wvalid[8 +: 1]),
    .AXI_08_WREADY(m_axi_hbm_int_wready[8 +: 1]),
    .AXI_08_BID(m_axi_hbm_int_bid[8*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_08_BRESP(m_axi_hbm_int_bresp[8*2 +: 2]),
    .AXI_08_BVALID(m_axi_hbm_int_bvalid[8 +: 1]),
    .AXI_08_BREADY(m_axi_hbm_int_bready[8 +: 1]),

    .AXI_09_ACLK(hbm_clk_int[9 +: 1]),
    .AXI_09_ARESET_N(!hbm_rst_int[9 +: 1]),

    .AXI_09_ARADDR(m_axi_hbm_int_araddr[9*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_09_ARBURST(m_axi_hbm_int_arburst[9*2 +: 2]),
    .AXI_09_ARID(m_axi_hbm_int_arid[9*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_09_ARLEN(m_axi_hbm_int_arlen[9*8 +: 4]),
    .AXI_09_ARSIZE(m_axi_hbm_int_arsize[9*3 +: 3]),
    .AXI_09_ARVALID(m_axi_hbm_int_arvalid[9 +: 1]),
    .AXI_09_ARREADY(m_axi_hbm_int_arready[9 +: 1]),
    .AXI_09_RDATA_PARITY(),
    .AXI_09_RDATA(m_axi_hbm_int_rdata[9*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_09_RID(m_axi_hbm_int_rid[9*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_09_RLAST(m_axi_hbm_int_rlast[9 +: 1]),
    .AXI_09_RRESP(m_axi_hbm_int_rresp[9*2 +: 2]),
    .AXI_09_RVALID(m_axi_hbm_int_rvalid[9 +: 1]),
    .AXI_09_RREADY(m_axi_hbm_int_rready[9 +: 1]),
    .AXI_09_AWADDR(m_axi_hbm_int_awaddr[9*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_09_AWBURST(m_axi_hbm_int_awburst[9*2 +: 2]),
    .AXI_09_AWID(m_axi_hbm_int_awid[9*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_09_AWLEN(m_axi_hbm_int_awlen[9*8 +: 4]),
    .AXI_09_AWSIZE(m_axi_hbm_int_awsize[9*3 +: 3]),
    .AXI_09_AWVALID(m_axi_hbm_int_awvalid[9 +: 1]),
    .AXI_09_AWREADY(m_axi_hbm_int_awready[9 +: 1]),
    .AXI_09_WDATA(m_axi_hbm_int_wdata[9*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_09_WLAST(m_axi_hbm_int_wlast[9 +: 1]),
    .AXI_09_WSTRB(m_axi_hbm_int_wstrb[9*AXI_HBM_STRB_WIDTH +: AXI_HBM_STRB_WIDTH]),
    .AXI_09_WDATA_PARITY(32'd0),
    .AXI_09_WVALID(m_axi_hbm_int_wvalid[9 +: 1]),
    .AXI_09_WREADY(m_axi_hbm_int_wready[9 +: 1]),
    .AXI_09_BID(m_axi_hbm_int_bid[9*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_09_BRESP(m_axi_hbm_int_bresp[9*2 +: 2]),
    .AXI_09_BVALID(m_axi_hbm_int_bvalid[9 +: 1]),
    .AXI_09_BREADY(m_axi_hbm_int_bready[9 +: 1]),

    .AXI_10_ACLK(hbm_clk_int[10 +: 1]),
    .AXI_10_ARESET_N(!hbm_rst_int[10 +: 1]),

    .AXI_10_ARADDR(m_axi_hbm_int_araddr[10*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_10_ARBURST(m_axi_hbm_int_arburst[10*2 +: 2]),
    .AXI_10_ARID(m_axi_hbm_int_arid[10*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_10_ARLEN(m_axi_hbm_int_arlen[10*8 +: 4]),
    .AXI_10_ARSIZE(m_axi_hbm_int_arsize[10*3 +: 3]),
    .AXI_10_ARVALID(m_axi_hbm_int_arvalid[10 +: 1]),
    .AXI_10_ARREADY(m_axi_hbm_int_arready[10 +: 1]),
    .AXI_10_RDATA_PARITY(),
    .AXI_10_RDATA(m_axi_hbm_int_rdata[10*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_10_RID(m_axi_hbm_int_rid[10*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_10_RLAST(m_axi_hbm_int_rlast[10 +: 1]),
    .AXI_10_RRESP(m_axi_hbm_int_rresp[10*2 +: 2]),
    .AXI_10_RVALID(m_axi_hbm_int_rvalid[10 +: 1]),
    .AXI_10_RREADY(m_axi_hbm_int_rready[10 +: 1]),
    .AXI_10_AWADDR(m_axi_hbm_int_awaddr[10*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_10_AWBURST(m_axi_hbm_int_awburst[10*2 +: 2]),
    .AXI_10_AWID(m_axi_hbm_int_awid[10*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_10_AWLEN(m_axi_hbm_int_awlen[10*8 +: 4]),
    .AXI_10_AWSIZE(m_axi_hbm_int_awsize[10*3 +: 3]),
    .AXI_10_AWVALID(m_axi_hbm_int_awvalid[10 +: 1]),
    .AXI_10_AWREADY(m_axi_hbm_int_awready[10 +: 1]),
    .AXI_10_WDATA(m_axi_hbm_int_wdata[10*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_10_WLAST(m_axi_hbm_int_wlast[10 +: 1]),
    .AXI_10_WSTRB(m_axi_hbm_int_wstrb[10*AXI_HBM_STRB_WIDTH +: AXI_HBM_STRB_WIDTH]),
    .AXI_10_WDATA_PARITY(32'd0),
    .AXI_10_WVALID(m_axi_hbm_int_wvalid[10 +: 1]),
    .AXI_10_WREADY(m_axi_hbm_int_wready[10 +: 1]),
    .AXI_10_BID(m_axi_hbm_int_bid[10*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_10_BRESP(m_axi_hbm_int_bresp[10*2 +: 2]),
    .AXI_10_BVALID(m_axi_hbm_int_bvalid[10 +: 1]),
    .AXI_10_BREADY(m_axi_hbm_int_bready[10 +: 1]),

    .AXI_11_ACLK(hbm_clk_int[11 +: 1]),
    .AXI_11_ARESET_N(!hbm_rst_int[11 +: 1]),

    .AXI_11_ARADDR(m_axi_hbm_int_araddr[11*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_11_ARBURST(m_axi_hbm_int_arburst[11*2 +: 2]),
    .AXI_11_ARID(m_axi_hbm_int_arid[11*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_11_ARLEN(m_axi_hbm_int_arlen[11*8 +: 4]),
    .AXI_11_ARSIZE(m_axi_hbm_int_arsize[11*3 +: 3]),
    .AXI_11_ARVALID(m_axi_hbm_int_arvalid[11 +: 1]),
    .AXI_11_ARREADY(m_axi_hbm_int_arready[11 +: 1]),
    .AXI_11_RDATA_PARITY(),
    .AXI_11_RDATA(m_axi_hbm_int_rdata[11*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_11_RID(m_axi_hbm_int_rid[11*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_11_RLAST(m_axi_hbm_int_rlast[11 +: 1]),
    .AXI_11_RRESP(m_axi_hbm_int_rresp[11*2 +: 2]),
    .AXI_11_RVALID(m_axi_hbm_int_rvalid[11 +: 1]),
    .AXI_11_RREADY(m_axi_hbm_int_rready[11 +: 1]),
    .AXI_11_AWADDR(m_axi_hbm_int_awaddr[11*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_11_AWBURST(m_axi_hbm_int_awburst[11*2 +: 2]),
    .AXI_11_AWID(m_axi_hbm_int_awid[11*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_11_AWLEN(m_axi_hbm_int_awlen[11*8 +: 4]),
    .AXI_11_AWSIZE(m_axi_hbm_int_awsize[11*3 +: 3]),
    .AXI_11_AWVALID(m_axi_hbm_int_awvalid[11 +: 1]),
    .AXI_11_AWREADY(m_axi_hbm_int_awready[11 +: 1]),
    .AXI_11_WDATA(m_axi_hbm_int_wdata[11*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_11_WLAST(m_axi_hbm_int_wlast[11 +: 1]),
    .AXI_11_WSTRB(m_axi_hbm_int_wstrb[11*AXI_HBM_STRB_WIDTH +: AXI_HBM_STRB_WIDTH]),
    .AXI_11_WDATA_PARITY(32'd0),
    .AXI_11_WVALID(m_axi_hbm_int_wvalid[11 +: 1]),
    .AXI_11_WREADY(m_axi_hbm_int_wready[11 +: 1]),
    .AXI_11_BID(m_axi_hbm_int_bid[11*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_11_BRESP(m_axi_hbm_int_bresp[11*2 +: 2]),
    .AXI_11_BVALID(m_axi_hbm_int_bvalid[11 +: 1]),
    .AXI_11_BREADY(m_axi_hbm_int_bready[11 +: 1]),

    .AXI_12_ACLK(hbm_clk_int[12 +: 1]),
    .AXI_12_ARESET_N(!hbm_rst_int[12 +: 1]),

    .AXI_12_ARADDR(m_axi_hbm_int_araddr[12*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_12_ARBURST(m_axi_hbm_int_arburst[12*2 +: 2]),
    .AXI_12_ARID(m_axi_hbm_int_arid[12*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_12_ARLEN(m_axi_hbm_int_arlen[12*8 +: 4]),
    .AXI_12_ARSIZE(m_axi_hbm_int_arsize[12*3 +: 3]),
    .AXI_12_ARVALID(m_axi_hbm_int_arvalid[12 +: 1]),
    .AXI_12_ARREADY(m_axi_hbm_int_arready[12 +: 1]),
    .AXI_12_RDATA_PARITY(),
    .AXI_12_RDATA(m_axi_hbm_int_rdata[12*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_12_RID(m_axi_hbm_int_rid[12*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_12_RLAST(m_axi_hbm_int_rlast[12 +: 1]),
    .AXI_12_RRESP(m_axi_hbm_int_rresp[12*2 +: 2]),
    .AXI_12_RVALID(m_axi_hbm_int_rvalid[12 +: 1]),
    .AXI_12_RREADY(m_axi_hbm_int_rready[12 +: 1]),
    .AXI_12_AWADDR(m_axi_hbm_int_awaddr[12*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_12_AWBURST(m_axi_hbm_int_awburst[12*2 +: 2]),
    .AXI_12_AWID(m_axi_hbm_int_awid[12*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_12_AWLEN(m_axi_hbm_int_awlen[12*8 +: 4]),
    .AXI_12_AWSIZE(m_axi_hbm_int_awsize[12*3 +: 3]),
    .AXI_12_AWVALID(m_axi_hbm_int_awvalid[12 +: 1]),
    .AXI_12_AWREADY(m_axi_hbm_int_awready[12 +: 1]),
    .AXI_12_WDATA(m_axi_hbm_int_wdata[12*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_12_WLAST(m_axi_hbm_int_wlast[12 +: 1]),
    .AXI_12_WSTRB(m_axi_hbm_int_wstrb[12*AXI_HBM_STRB_WIDTH +: AXI_HBM_STRB_WIDTH]),
    .AXI_12_WDATA_PARITY(32'd0),
    .AXI_12_WVALID(m_axi_hbm_int_wvalid[12 +: 1]),
    .AXI_12_WREADY(m_axi_hbm_int_wready[12 +: 1]),
    .AXI_12_BID(m_axi_hbm_int_bid[12*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_12_BRESP(m_axi_hbm_int_bresp[12*2 +: 2]),
    .AXI_12_BVALID(m_axi_hbm_int_bvalid[12 +: 1]),
    .AXI_12_BREADY(m_axi_hbm_int_bready[12 +: 1]),

    .AXI_13_ACLK(hbm_clk_int[13 +: 1]),
    .AXI_13_ARESET_N(!hbm_rst_int[13 +: 1]),

    .AXI_13_ARADDR(m_axi_hbm_int_araddr[13*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_13_ARBURST(m_axi_hbm_int_arburst[13*2 +: 2]),
    .AXI_13_ARID(m_axi_hbm_int_arid[13*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_13_ARLEN(m_axi_hbm_int_arlen[13*8 +: 4]),
    .AXI_13_ARSIZE(m_axi_hbm_int_arsize[13*3 +: 3]),
    .AXI_13_ARVALID(m_axi_hbm_int_arvalid[13 +: 1]),
    .AXI_13_ARREADY(m_axi_hbm_int_arready[13 +: 1]),
    .AXI_13_RDATA_PARITY(),
    .AXI_13_RDATA(m_axi_hbm_int_rdata[13*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_13_RID(m_axi_hbm_int_rid[13*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_13_RLAST(m_axi_hbm_int_rlast[13 +: 1]),
    .AXI_13_RRESP(m_axi_hbm_int_rresp[13*2 +: 2]),
    .AXI_13_RVALID(m_axi_hbm_int_rvalid[13 +: 1]),
    .AXI_13_RREADY(m_axi_hbm_int_rready[13 +: 1]),
    .AXI_13_AWADDR(m_axi_hbm_int_awaddr[13*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_13_AWBURST(m_axi_hbm_int_awburst[13*2 +: 2]),
    .AXI_13_AWID(m_axi_hbm_int_awid[13*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_13_AWLEN(m_axi_hbm_int_awlen[13*8 +: 4]),
    .AXI_13_AWSIZE(m_axi_hbm_int_awsize[13*3 +: 3]),
    .AXI_13_AWVALID(m_axi_hbm_int_awvalid[13 +: 1]),
    .AXI_13_AWREADY(m_axi_hbm_int_awready[13 +: 1]),
    .AXI_13_WDATA(m_axi_hbm_int_wdata[13*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_13_WLAST(m_axi_hbm_int_wlast[13 +: 1]),
    .AXI_13_WSTRB(m_axi_hbm_int_wstrb[13*AXI_HBM_STRB_WIDTH +: AXI_HBM_STRB_WIDTH]),
    .AXI_13_WDATA_PARITY(32'd0),
    .AXI_13_WVALID(m_axi_hbm_int_wvalid[13 +: 1]),
    .AXI_13_WREADY(m_axi_hbm_int_wready[13 +: 1]),
    .AXI_13_BID(m_axi_hbm_int_bid[13*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_13_BRESP(m_axi_hbm_int_bresp[13*2 +: 2]),
    .AXI_13_BVALID(m_axi_hbm_int_bvalid[13 +: 1]),
    .AXI_13_BREADY(m_axi_hbm_int_bready[13 +: 1]),

    .AXI_14_ACLK(hbm_clk_int[14 +: 1]),
    .AXI_14_ARESET_N(!hbm_rst_int[14 +: 1]),

    .AXI_14_ARADDR(m_axi_hbm_int_araddr[14*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_14_ARBURST(m_axi_hbm_int_arburst[14*2 +: 2]),
    .AXI_14_ARID(m_axi_hbm_int_arid[14*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_14_ARLEN(m_axi_hbm_int_arlen[14*8 +: 4]),
    .AXI_14_ARSIZE(m_axi_hbm_int_arsize[14*3 +: 3]),
    .AXI_14_ARVALID(m_axi_hbm_int_arvalid[14 +: 1]),
    .AXI_14_ARREADY(m_axi_hbm_int_arready[14 +: 1]),
    .AXI_14_RDATA_PARITY(),
    .AXI_14_RDATA(m_axi_hbm_int_rdata[14*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_14_RID(m_axi_hbm_int_rid[14*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_14_RLAST(m_axi_hbm_int_rlast[14 +: 1]),
    .AXI_14_RRESP(m_axi_hbm_int_rresp[14*2 +: 2]),
    .AXI_14_RVALID(m_axi_hbm_int_rvalid[14 +: 1]),
    .AXI_14_RREADY(m_axi_hbm_int_rready[14 +: 1]),
    .AXI_14_AWADDR(m_axi_hbm_int_awaddr[14*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_14_AWBURST(m_axi_hbm_int_awburst[14*2 +: 2]),
    .AXI_14_AWID(m_axi_hbm_int_awid[14*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_14_AWLEN(m_axi_hbm_int_awlen[14*8 +: 4]),
    .AXI_14_AWSIZE(m_axi_hbm_int_awsize[14*3 +: 3]),
    .AXI_14_AWVALID(m_axi_hbm_int_awvalid[14 +: 1]),
    .AXI_14_AWREADY(m_axi_hbm_int_awready[14 +: 1]),
    .AXI_14_WDATA(m_axi_hbm_int_wdata[14*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_14_WLAST(m_axi_hbm_int_wlast[14 +: 1]),
    .AXI_14_WSTRB(m_axi_hbm_int_wstrb[14*AXI_HBM_STRB_WIDTH +: AXI_HBM_STRB_WIDTH]),
    .AXI_14_WDATA_PARITY(32'd0),
    .AXI_14_WVALID(m_axi_hbm_int_wvalid[14 +: 1]),
    .AXI_14_WREADY(m_axi_hbm_int_wready[14 +: 1]),
    .AXI_14_BID(m_axi_hbm_int_bid[14*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_14_BRESP(m_axi_hbm_int_bresp[14*2 +: 2]),
    .AXI_14_BVALID(m_axi_hbm_int_bvalid[14 +: 1]),
    .AXI_14_BREADY(m_axi_hbm_int_bready[14 +: 1]),

    .AXI_15_ACLK(hbm_clk_int[15 +: 1]),
    .AXI_15_ARESET_N(!hbm_rst_int[15 +: 1]),

    .AXI_15_ARADDR(m_axi_hbm_int_araddr[15*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_15_ARBURST(m_axi_hbm_int_arburst[15*2 +: 2]),
    .AXI_15_ARID(m_axi_hbm_int_arid[15*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_15_ARLEN(m_axi_hbm_int_arlen[15*8 +: 4]),
    .AXI_15_ARSIZE(m_axi_hbm_int_arsize[15*3 +: 3]),
    .AXI_15_ARVALID(m_axi_hbm_int_arvalid[15 +: 1]),
    .AXI_15_ARREADY(m_axi_hbm_int_arready[15 +: 1]),
    .AXI_15_RDATA_PARITY(),
    .AXI_15_RDATA(m_axi_hbm_int_rdata[15*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_15_RID(m_axi_hbm_int_rid[15*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_15_RLAST(m_axi_hbm_int_rlast[15 +: 1]),
    .AXI_15_RRESP(m_axi_hbm_int_rresp[15*2 +: 2]),
    .AXI_15_RVALID(m_axi_hbm_int_rvalid[15 +: 1]),
    .AXI_15_RREADY(m_axi_hbm_int_rready[15 +: 1]),
    .AXI_15_AWADDR(m_axi_hbm_int_awaddr[15*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_15_AWBURST(m_axi_hbm_int_awburst[15*2 +: 2]),
    .AXI_15_AWID(m_axi_hbm_int_awid[15*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_15_AWLEN(m_axi_hbm_int_awlen[15*8 +: 4]),
    .AXI_15_AWSIZE(m_axi_hbm_int_awsize[15*3 +: 3]),
    .AXI_15_AWVALID(m_axi_hbm_int_awvalid[15 +: 1]),
    .AXI_15_AWREADY(m_axi_hbm_int_awready[15 +: 1]),
    .AXI_15_WDATA(m_axi_hbm_int_wdata[15*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_15_WLAST(m_axi_hbm_int_wlast[15 +: 1]),
    .AXI_15_WSTRB(m_axi_hbm_int_wstrb[15*AXI_HBM_STRB_WIDTH +: AXI_HBM_STRB_WIDTH]),
    .AXI_15_WDATA_PARITY(32'd0),
    .AXI_15_WVALID(m_axi_hbm_int_wvalid[15 +: 1]),
    .AXI_15_WREADY(m_axi_hbm_int_wready[15 +: 1]),
    .AXI_15_BID(m_axi_hbm_int_bid[15*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_15_BRESP(m_axi_hbm_int_bresp[15*2 +: 2]),
    .AXI_15_BVALID(m_axi_hbm_int_bvalid[15 +: 1]),
    .AXI_15_BREADY(m_axi_hbm_int_bready[15 +: 1]),

    .AXI_16_ACLK(hbm_clk_int[16 +: 1]),
    .AXI_16_ARESET_N(!hbm_rst_int[16 +: 1]),

    .AXI_16_ARADDR(m_axi_hbm_int_araddr[16*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_16_ARBURST(m_axi_hbm_int_arburst[16*2 +: 2]),
    .AXI_16_ARID(m_axi_hbm_int_arid[16*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_16_ARLEN(m_axi_hbm_int_arlen[16*8 +: 4]),
    .AXI_16_ARSIZE(m_axi_hbm_int_arsize[16*3 +: 3]),
    .AXI_16_ARVALID(m_axi_hbm_int_arvalid[16 +: 1]),
    .AXI_16_ARREADY(m_axi_hbm_int_arready[16 +: 1]),
    .AXI_16_RDATA_PARITY(),
    .AXI_16_RDATA(m_axi_hbm_int_rdata[16*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_16_RID(m_axi_hbm_int_rid[16*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_16_RLAST(m_axi_hbm_int_rlast[16 +: 1]),
    .AXI_16_RRESP(m_axi_hbm_int_rresp[16*2 +: 2]),
    .AXI_16_RVALID(m_axi_hbm_int_rvalid[16 +: 1]),
    .AXI_16_RREADY(m_axi_hbm_int_rready[16 +: 1]),
    .AXI_16_AWADDR(m_axi_hbm_int_awaddr[16*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_16_AWBURST(m_axi_hbm_int_awburst[16*2 +: 2]),
    .AXI_16_AWID(m_axi_hbm_int_awid[16*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_16_AWLEN(m_axi_hbm_int_awlen[16*8 +: 4]),
    .AXI_16_AWSIZE(m_axi_hbm_int_awsize[16*3 +: 3]),
    .AXI_16_AWVALID(m_axi_hbm_int_awvalid[16 +: 1]),
    .AXI_16_AWREADY(m_axi_hbm_int_awready[16 +: 1]),
    .AXI_16_WDATA(m_axi_hbm_int_wdata[16*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_16_WLAST(m_axi_hbm_int_wlast[16 +: 1]),
    .AXI_16_WSTRB(m_axi_hbm_int_wstrb[16*AXI_HBM_STRB_WIDTH +: AXI_HBM_STRB_WIDTH]),
    .AXI_16_WDATA_PARITY(32'd0),
    .AXI_16_WVALID(m_axi_hbm_int_wvalid[16 +: 1]),
    .AXI_16_WREADY(m_axi_hbm_int_wready[16 +: 1]),
    .AXI_16_BID(m_axi_hbm_int_bid[16*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_16_BRESP(m_axi_hbm_int_bresp[16*2 +: 2]),
    .AXI_16_BVALID(m_axi_hbm_int_bvalid[16 +: 1]),
    .AXI_16_BREADY(m_axi_hbm_int_bready[16 +: 1]),

    .AXI_17_ACLK(hbm_clk_int[17 +: 1]),
    .AXI_17_ARESET_N(!hbm_rst_int[17 +: 1]),

    .AXI_17_ARADDR(m_axi_hbm_int_araddr[17*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_17_ARBURST(m_axi_hbm_int_arburst[17*2 +: 2]),
    .AXI_17_ARID(m_axi_hbm_int_arid[17*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_17_ARLEN(m_axi_hbm_int_arlen[17*8 +: 4]),
    .AXI_17_ARSIZE(m_axi_hbm_int_arsize[17*3 +: 3]),
    .AXI_17_ARVALID(m_axi_hbm_int_arvalid[17 +: 1]),
    .AXI_17_ARREADY(m_axi_hbm_int_arready[17 +: 1]),
    .AXI_17_RDATA_PARITY(),
    .AXI_17_RDATA(m_axi_hbm_int_rdata[17*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_17_RID(m_axi_hbm_int_rid[17*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_17_RLAST(m_axi_hbm_int_rlast[17 +: 1]),
    .AXI_17_RRESP(m_axi_hbm_int_rresp[17*2 +: 2]),
    .AXI_17_RVALID(m_axi_hbm_int_rvalid[17 +: 1]),
    .AXI_17_RREADY(m_axi_hbm_int_rready[17 +: 1]),
    .AXI_17_AWADDR(m_axi_hbm_int_awaddr[17*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_17_AWBURST(m_axi_hbm_int_awburst[17*2 +: 2]),
    .AXI_17_AWID(m_axi_hbm_int_awid[17*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_17_AWLEN(m_axi_hbm_int_awlen[17*8 +: 4]),
    .AXI_17_AWSIZE(m_axi_hbm_int_awsize[17*3 +: 3]),
    .AXI_17_AWVALID(m_axi_hbm_int_awvalid[17 +: 1]),
    .AXI_17_AWREADY(m_axi_hbm_int_awready[17 +: 1]),
    .AXI_17_WDATA(m_axi_hbm_int_wdata[17*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_17_WLAST(m_axi_hbm_int_wlast[17 +: 1]),
    .AXI_17_WSTRB(m_axi_hbm_int_wstrb[17*AXI_HBM_STRB_WIDTH +: AXI_HBM_STRB_WIDTH]),
    .AXI_17_WDATA_PARITY(32'd0),
    .AXI_17_WVALID(m_axi_hbm_int_wvalid[17 +: 1]),
    .AXI_17_WREADY(m_axi_hbm_int_wready[17 +: 1]),
    .AXI_17_BID(m_axi_hbm_int_bid[17*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_17_BRESP(m_axi_hbm_int_bresp[17*2 +: 2]),
    .AXI_17_BVALID(m_axi_hbm_int_bvalid[17 +: 1]),
    .AXI_17_BREADY(m_axi_hbm_int_bready[17 +: 1]),

    .AXI_18_ACLK(hbm_clk_int[18 +: 1]),
    .AXI_18_ARESET_N(!hbm_rst_int[18 +: 1]),

    .AXI_18_ARADDR(m_axi_hbm_int_araddr[18*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_18_ARBURST(m_axi_hbm_int_arburst[18*2 +: 2]),
    .AXI_18_ARID(m_axi_hbm_int_arid[18*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_18_ARLEN(m_axi_hbm_int_arlen[18*8 +: 4]),
    .AXI_18_ARSIZE(m_axi_hbm_int_arsize[18*3 +: 3]),
    .AXI_18_ARVALID(m_axi_hbm_int_arvalid[18 +: 1]),
    .AXI_18_ARREADY(m_axi_hbm_int_arready[18 +: 1]),
    .AXI_18_RDATA_PARITY(),
    .AXI_18_RDATA(m_axi_hbm_int_rdata[18*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_18_RID(m_axi_hbm_int_rid[18*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_18_RLAST(m_axi_hbm_int_rlast[18 +: 1]),
    .AXI_18_RRESP(m_axi_hbm_int_rresp[18*2 +: 2]),
    .AXI_18_RVALID(m_axi_hbm_int_rvalid[18 +: 1]),
    .AXI_18_RREADY(m_axi_hbm_int_rready[18 +: 1]),
    .AXI_18_AWADDR(m_axi_hbm_int_awaddr[18*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_18_AWBURST(m_axi_hbm_int_awburst[18*2 +: 2]),
    .AXI_18_AWID(m_axi_hbm_int_awid[18*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_18_AWLEN(m_axi_hbm_int_awlen[18*8 +: 4]),
    .AXI_18_AWSIZE(m_axi_hbm_int_awsize[18*3 +: 3]),
    .AXI_18_AWVALID(m_axi_hbm_int_awvalid[18 +: 1]),
    .AXI_18_AWREADY(m_axi_hbm_int_awready[18 +: 1]),
    .AXI_18_WDATA(m_axi_hbm_int_wdata[18*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_18_WLAST(m_axi_hbm_int_wlast[18 +: 1]),
    .AXI_18_WSTRB(m_axi_hbm_int_wstrb[18*AXI_HBM_STRB_WIDTH +: AXI_HBM_STRB_WIDTH]),
    .AXI_18_WDATA_PARITY(32'd0),
    .AXI_18_WVALID(m_axi_hbm_int_wvalid[18 +: 1]),
    .AXI_18_WREADY(m_axi_hbm_int_wready[18 +: 1]),
    .AXI_18_BID(m_axi_hbm_int_bid[18*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_18_BRESP(m_axi_hbm_int_bresp[18*2 +: 2]),
    .AXI_18_BVALID(m_axi_hbm_int_bvalid[18 +: 1]),
    .AXI_18_BREADY(m_axi_hbm_int_bready[18 +: 1]),

    .AXI_19_ACLK(hbm_clk_int[19 +: 1]),
    .AXI_19_ARESET_N(!hbm_rst_int[19 +: 1]),

    .AXI_19_ARADDR(m_axi_hbm_int_araddr[19*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_19_ARBURST(m_axi_hbm_int_arburst[19*2 +: 2]),
    .AXI_19_ARID(m_axi_hbm_int_arid[19*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_19_ARLEN(m_axi_hbm_int_arlen[19*8 +: 4]),
    .AXI_19_ARSIZE(m_axi_hbm_int_arsize[19*3 +: 3]),
    .AXI_19_ARVALID(m_axi_hbm_int_arvalid[19 +: 1]),
    .AXI_19_ARREADY(m_axi_hbm_int_arready[19 +: 1]),
    .AXI_19_RDATA_PARITY(),
    .AXI_19_RDATA(m_axi_hbm_int_rdata[19*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_19_RID(m_axi_hbm_int_rid[19*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_19_RLAST(m_axi_hbm_int_rlast[19 +: 1]),
    .AXI_19_RRESP(m_axi_hbm_int_rresp[19*2 +: 2]),
    .AXI_19_RVALID(m_axi_hbm_int_rvalid[19 +: 1]),
    .AXI_19_RREADY(m_axi_hbm_int_rready[19 +: 1]),
    .AXI_19_AWADDR(m_axi_hbm_int_awaddr[19*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_19_AWBURST(m_axi_hbm_int_awburst[19*2 +: 2]),
    .AXI_19_AWID(m_axi_hbm_int_awid[19*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_19_AWLEN(m_axi_hbm_int_awlen[19*8 +: 4]),
    .AXI_19_AWSIZE(m_axi_hbm_int_awsize[19*3 +: 3]),
    .AXI_19_AWVALID(m_axi_hbm_int_awvalid[19 +: 1]),
    .AXI_19_AWREADY(m_axi_hbm_int_awready[19 +: 1]),
    .AXI_19_WDATA(m_axi_hbm_int_wdata[19*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_19_WLAST(m_axi_hbm_int_wlast[19 +: 1]),
    .AXI_19_WSTRB(m_axi_hbm_int_wstrb[19*AXI_HBM_STRB_WIDTH +: AXI_HBM_STRB_WIDTH]),
    .AXI_19_WDATA_PARITY(32'd0),
    .AXI_19_WVALID(m_axi_hbm_int_wvalid[19 +: 1]),
    .AXI_19_WREADY(m_axi_hbm_int_wready[19 +: 1]),
    .AXI_19_BID(m_axi_hbm_int_bid[19*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_19_BRESP(m_axi_hbm_int_bresp[19*2 +: 2]),
    .AXI_19_BVALID(m_axi_hbm_int_bvalid[19 +: 1]),
    .AXI_19_BREADY(m_axi_hbm_int_bready[19 +: 1]),

    .AXI_20_ACLK(hbm_clk_int[20 +: 1]),
    .AXI_20_ARESET_N(!hbm_rst_int[20 +: 1]),

    .AXI_20_ARADDR(m_axi_hbm_int_araddr[20*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_20_ARBURST(m_axi_hbm_int_arburst[20*2 +: 2]),
    .AXI_20_ARID(m_axi_hbm_int_arid[20*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_20_ARLEN(m_axi_hbm_int_arlen[20*8 +: 4]),
    .AXI_20_ARSIZE(m_axi_hbm_int_arsize[20*3 +: 3]),
    .AXI_20_ARVALID(m_axi_hbm_int_arvalid[20 +: 1]),
    .AXI_20_ARREADY(m_axi_hbm_int_arready[20 +: 1]),
    .AXI_20_RDATA_PARITY(),
    .AXI_20_RDATA(m_axi_hbm_int_rdata[20*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_20_RID(m_axi_hbm_int_rid[20*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_20_RLAST(m_axi_hbm_int_rlast[20 +: 1]),
    .AXI_20_RRESP(m_axi_hbm_int_rresp[20*2 +: 2]),
    .AXI_20_RVALID(m_axi_hbm_int_rvalid[20 +: 1]),
    .AXI_20_RREADY(m_axi_hbm_int_rready[20 +: 1]),
    .AXI_20_AWADDR(m_axi_hbm_int_awaddr[20*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_20_AWBURST(m_axi_hbm_int_awburst[20*2 +: 2]),
    .AXI_20_AWID(m_axi_hbm_int_awid[20*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_20_AWLEN(m_axi_hbm_int_awlen[20*8 +: 4]),
    .AXI_20_AWSIZE(m_axi_hbm_int_awsize[20*3 +: 3]),
    .AXI_20_AWVALID(m_axi_hbm_int_awvalid[20 +: 1]),
    .AXI_20_AWREADY(m_axi_hbm_int_awready[20 +: 1]),
    .AXI_20_WDATA(m_axi_hbm_int_wdata[20*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_20_WLAST(m_axi_hbm_int_wlast[20 +: 1]),
    .AXI_20_WSTRB(m_axi_hbm_int_wstrb[20*AXI_HBM_STRB_WIDTH +: AXI_HBM_STRB_WIDTH]),
    .AXI_20_WDATA_PARITY(32'd0),
    .AXI_20_WVALID(m_axi_hbm_int_wvalid[20 +: 1]),
    .AXI_20_WREADY(m_axi_hbm_int_wready[20 +: 1]),
    .AXI_20_BID(m_axi_hbm_int_bid[20*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_20_BRESP(m_axi_hbm_int_bresp[20*2 +: 2]),
    .AXI_20_BVALID(m_axi_hbm_int_bvalid[20 +: 1]),
    .AXI_20_BREADY(m_axi_hbm_int_bready[20 +: 1]),

    .AXI_21_ACLK(hbm_clk_int[21 +: 1]),
    .AXI_21_ARESET_N(!hbm_rst_int[21 +: 1]),

    .AXI_21_ARADDR(m_axi_hbm_int_araddr[21*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_21_ARBURST(m_axi_hbm_int_arburst[21*2 +: 2]),
    .AXI_21_ARID(m_axi_hbm_int_arid[21*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_21_ARLEN(m_axi_hbm_int_arlen[21*8 +: 4]),
    .AXI_21_ARSIZE(m_axi_hbm_int_arsize[21*3 +: 3]),
    .AXI_21_ARVALID(m_axi_hbm_int_arvalid[21 +: 1]),
    .AXI_21_ARREADY(m_axi_hbm_int_arready[21 +: 1]),
    .AXI_21_RDATA_PARITY(),
    .AXI_21_RDATA(m_axi_hbm_int_rdata[21*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_21_RID(m_axi_hbm_int_rid[21*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_21_RLAST(m_axi_hbm_int_rlast[21 +: 1]),
    .AXI_21_RRESP(m_axi_hbm_int_rresp[21*2 +: 2]),
    .AXI_21_RVALID(m_axi_hbm_int_rvalid[21 +: 1]),
    .AXI_21_RREADY(m_axi_hbm_int_rready[21 +: 1]),
    .AXI_21_AWADDR(m_axi_hbm_int_awaddr[21*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_21_AWBURST(m_axi_hbm_int_awburst[21*2 +: 2]),
    .AXI_21_AWID(m_axi_hbm_int_awid[21*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_21_AWLEN(m_axi_hbm_int_awlen[21*8 +: 4]),
    .AXI_21_AWSIZE(m_axi_hbm_int_awsize[21*3 +: 3]),
    .AXI_21_AWVALID(m_axi_hbm_int_awvalid[21 +: 1]),
    .AXI_21_AWREADY(m_axi_hbm_int_awready[21 +: 1]),
    .AXI_21_WDATA(m_axi_hbm_int_wdata[21*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_21_WLAST(m_axi_hbm_int_wlast[21 +: 1]),
    .AXI_21_WSTRB(m_axi_hbm_int_wstrb[21*AXI_HBM_STRB_WIDTH +: AXI_HBM_STRB_WIDTH]),
    .AXI_21_WDATA_PARITY(32'd0),
    .AXI_21_WVALID(m_axi_hbm_int_wvalid[21 +: 1]),
    .AXI_21_WREADY(m_axi_hbm_int_wready[21 +: 1]),
    .AXI_21_BID(m_axi_hbm_int_bid[21*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_21_BRESP(m_axi_hbm_int_bresp[21*2 +: 2]),
    .AXI_21_BVALID(m_axi_hbm_int_bvalid[21 +: 1]),
    .AXI_21_BREADY(m_axi_hbm_int_bready[21 +: 1]),

    .AXI_22_ACLK(hbm_clk_int[22 +: 1]),
    .AXI_22_ARESET_N(!hbm_rst_int[22 +: 1]),

    .AXI_22_ARADDR(m_axi_hbm_int_araddr[22*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_22_ARBURST(m_axi_hbm_int_arburst[22*2 +: 2]),
    .AXI_22_ARID(m_axi_hbm_int_arid[22*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_22_ARLEN(m_axi_hbm_int_arlen[22*8 +: 4]),
    .AXI_22_ARSIZE(m_axi_hbm_int_arsize[22*3 +: 3]),
    .AXI_22_ARVALID(m_axi_hbm_int_arvalid[22 +: 1]),
    .AXI_22_ARREADY(m_axi_hbm_int_arready[22 +: 1]),
    .AXI_22_RDATA_PARITY(),
    .AXI_22_RDATA(m_axi_hbm_int_rdata[22*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_22_RID(m_axi_hbm_int_rid[22*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_22_RLAST(m_axi_hbm_int_rlast[22 +: 1]),
    .AXI_22_RRESP(m_axi_hbm_int_rresp[22*2 +: 2]),
    .AXI_22_RVALID(m_axi_hbm_int_rvalid[22 +: 1]),
    .AXI_22_RREADY(m_axi_hbm_int_rready[22 +: 1]),
    .AXI_22_AWADDR(m_axi_hbm_int_awaddr[22*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_22_AWBURST(m_axi_hbm_int_awburst[22*2 +: 2]),
    .AXI_22_AWID(m_axi_hbm_int_awid[22*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_22_AWLEN(m_axi_hbm_int_awlen[22*8 +: 4]),
    .AXI_22_AWSIZE(m_axi_hbm_int_awsize[22*3 +: 3]),
    .AXI_22_AWVALID(m_axi_hbm_int_awvalid[22 +: 1]),
    .AXI_22_AWREADY(m_axi_hbm_int_awready[22 +: 1]),
    .AXI_22_WDATA(m_axi_hbm_int_wdata[22*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_22_WLAST(m_axi_hbm_int_wlast[22 +: 1]),
    .AXI_22_WSTRB(m_axi_hbm_int_wstrb[22*AXI_HBM_STRB_WIDTH +: AXI_HBM_STRB_WIDTH]),
    .AXI_22_WDATA_PARITY(32'd0),
    .AXI_22_WVALID(m_axi_hbm_int_wvalid[22 +: 1]),
    .AXI_22_WREADY(m_axi_hbm_int_wready[22 +: 1]),
    .AXI_22_BID(m_axi_hbm_int_bid[22*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_22_BRESP(m_axi_hbm_int_bresp[22*2 +: 2]),
    .AXI_22_BVALID(m_axi_hbm_int_bvalid[22 +: 1]),
    .AXI_22_BREADY(m_axi_hbm_int_bready[22 +: 1]),

    .AXI_23_ACLK(hbm_clk_int[23 +: 1]),
    .AXI_23_ARESET_N(!hbm_rst_int[23 +: 1]),

    .AXI_23_ARADDR(m_axi_hbm_int_araddr[23*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_23_ARBURST(m_axi_hbm_int_arburst[23*2 +: 2]),
    .AXI_23_ARID(m_axi_hbm_int_arid[23*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_23_ARLEN(m_axi_hbm_int_arlen[23*8 +: 4]),
    .AXI_23_ARSIZE(m_axi_hbm_int_arsize[23*3 +: 3]),
    .AXI_23_ARVALID(m_axi_hbm_int_arvalid[23 +: 1]),
    .AXI_23_ARREADY(m_axi_hbm_int_arready[23 +: 1]),
    .AXI_23_RDATA_PARITY(),
    .AXI_23_RDATA(m_axi_hbm_int_rdata[23*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_23_RID(m_axi_hbm_int_rid[23*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_23_RLAST(m_axi_hbm_int_rlast[23 +: 1]),
    .AXI_23_RRESP(m_axi_hbm_int_rresp[23*2 +: 2]),
    .AXI_23_RVALID(m_axi_hbm_int_rvalid[23 +: 1]),
    .AXI_23_RREADY(m_axi_hbm_int_rready[23 +: 1]),
    .AXI_23_AWADDR(m_axi_hbm_int_awaddr[23*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_23_AWBURST(m_axi_hbm_int_awburst[23*2 +: 2]),
    .AXI_23_AWID(m_axi_hbm_int_awid[23*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_23_AWLEN(m_axi_hbm_int_awlen[23*8 +: 4]),
    .AXI_23_AWSIZE(m_axi_hbm_int_awsize[23*3 +: 3]),
    .AXI_23_AWVALID(m_axi_hbm_int_awvalid[23 +: 1]),
    .AXI_23_AWREADY(m_axi_hbm_int_awready[23 +: 1]),
    .AXI_23_WDATA(m_axi_hbm_int_wdata[23*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_23_WLAST(m_axi_hbm_int_wlast[23 +: 1]),
    .AXI_23_WSTRB(m_axi_hbm_int_wstrb[23*AXI_HBM_STRB_WIDTH +: AXI_HBM_STRB_WIDTH]),
    .AXI_23_WDATA_PARITY(32'd0),
    .AXI_23_WVALID(m_axi_hbm_int_wvalid[23 +: 1]),
    .AXI_23_WREADY(m_axi_hbm_int_wready[23 +: 1]),
    .AXI_23_BID(m_axi_hbm_int_bid[23*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_23_BRESP(m_axi_hbm_int_bresp[23*2 +: 2]),
    .AXI_23_BVALID(m_axi_hbm_int_bvalid[23 +: 1]),
    .AXI_23_BREADY(m_axi_hbm_int_bready[23 +: 1]),

    .AXI_24_ACLK(hbm_clk_int[24 +: 1]),
    .AXI_24_ARESET_N(!hbm_rst_int[24 +: 1]),

    .AXI_24_ARADDR(m_axi_hbm_int_araddr[24*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_24_ARBURST(m_axi_hbm_int_arburst[24*2 +: 2]),
    .AXI_24_ARID(m_axi_hbm_int_arid[24*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_24_ARLEN(m_axi_hbm_int_arlen[24*8 +: 4]),
    .AXI_24_ARSIZE(m_axi_hbm_int_arsize[24*3 +: 3]),
    .AXI_24_ARVALID(m_axi_hbm_int_arvalid[24 +: 1]),
    .AXI_24_ARREADY(m_axi_hbm_int_arready[24 +: 1]),
    .AXI_24_RDATA_PARITY(),
    .AXI_24_RDATA(m_axi_hbm_int_rdata[24*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_24_RID(m_axi_hbm_int_rid[24*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_24_RLAST(m_axi_hbm_int_rlast[24 +: 1]),
    .AXI_24_RRESP(m_axi_hbm_int_rresp[24*2 +: 2]),
    .AXI_24_RVALID(m_axi_hbm_int_rvalid[24 +: 1]),
    .AXI_24_RREADY(m_axi_hbm_int_rready[24 +: 1]),
    .AXI_24_AWADDR(m_axi_hbm_int_awaddr[24*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_24_AWBURST(m_axi_hbm_int_awburst[24*2 +: 2]),
    .AXI_24_AWID(m_axi_hbm_int_awid[24*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_24_AWLEN(m_axi_hbm_int_awlen[24*8 +: 4]),
    .AXI_24_AWSIZE(m_axi_hbm_int_awsize[24*3 +: 3]),
    .AXI_24_AWVALID(m_axi_hbm_int_awvalid[24 +: 1]),
    .AXI_24_AWREADY(m_axi_hbm_int_awready[24 +: 1]),
    .AXI_24_WDATA(m_axi_hbm_int_wdata[24*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_24_WLAST(m_axi_hbm_int_wlast[24 +: 1]),
    .AXI_24_WSTRB(m_axi_hbm_int_wstrb[24*AXI_HBM_STRB_WIDTH +: AXI_HBM_STRB_WIDTH]),
    .AXI_24_WDATA_PARITY(32'd0),
    .AXI_24_WVALID(m_axi_hbm_int_wvalid[24 +: 1]),
    .AXI_24_WREADY(m_axi_hbm_int_wready[24 +: 1]),
    .AXI_24_BID(m_axi_hbm_int_bid[24*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_24_BRESP(m_axi_hbm_int_bresp[24*2 +: 2]),
    .AXI_24_BVALID(m_axi_hbm_int_bvalid[24 +: 1]),
    .AXI_24_BREADY(m_axi_hbm_int_bready[24 +: 1]),

    .AXI_25_ACLK(hbm_clk_int[25 +: 1]),
    .AXI_25_ARESET_N(!hbm_rst_int[25 +: 1]),

    .AXI_25_ARADDR(m_axi_hbm_int_araddr[25*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_25_ARBURST(m_axi_hbm_int_arburst[25*2 +: 2]),
    .AXI_25_ARID(m_axi_hbm_int_arid[25*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_25_ARLEN(m_axi_hbm_int_arlen[25*8 +: 4]),
    .AXI_25_ARSIZE(m_axi_hbm_int_arsize[25*3 +: 3]),
    .AXI_25_ARVALID(m_axi_hbm_int_arvalid[25 +: 1]),
    .AXI_25_ARREADY(m_axi_hbm_int_arready[25 +: 1]),
    .AXI_25_RDATA_PARITY(),
    .AXI_25_RDATA(m_axi_hbm_int_rdata[25*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_25_RID(m_axi_hbm_int_rid[25*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_25_RLAST(m_axi_hbm_int_rlast[25 +: 1]),
    .AXI_25_RRESP(m_axi_hbm_int_rresp[25*2 +: 2]),
    .AXI_25_RVALID(m_axi_hbm_int_rvalid[25 +: 1]),
    .AXI_25_RREADY(m_axi_hbm_int_rready[25 +: 1]),
    .AXI_25_AWADDR(m_axi_hbm_int_awaddr[25*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_25_AWBURST(m_axi_hbm_int_awburst[25*2 +: 2]),
    .AXI_25_AWID(m_axi_hbm_int_awid[25*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_25_AWLEN(m_axi_hbm_int_awlen[25*8 +: 4]),
    .AXI_25_AWSIZE(m_axi_hbm_int_awsize[25*3 +: 3]),
    .AXI_25_AWVALID(m_axi_hbm_int_awvalid[25 +: 1]),
    .AXI_25_AWREADY(m_axi_hbm_int_awready[25 +: 1]),
    .AXI_25_WDATA(m_axi_hbm_int_wdata[25*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_25_WLAST(m_axi_hbm_int_wlast[25 +: 1]),
    .AXI_25_WSTRB(m_axi_hbm_int_wstrb[25*AXI_HBM_STRB_WIDTH +: AXI_HBM_STRB_WIDTH]),
    .AXI_25_WDATA_PARITY(32'd0),
    .AXI_25_WVALID(m_axi_hbm_int_wvalid[25 +: 1]),
    .AXI_25_WREADY(m_axi_hbm_int_wready[25 +: 1]),
    .AXI_25_BID(m_axi_hbm_int_bid[25*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_25_BRESP(m_axi_hbm_int_bresp[25*2 +: 2]),
    .AXI_25_BVALID(m_axi_hbm_int_bvalid[25 +: 1]),
    .AXI_25_BREADY(m_axi_hbm_int_bready[25 +: 1]),

    .AXI_26_ACLK(hbm_clk_int[26 +: 1]),
    .AXI_26_ARESET_N(!hbm_rst_int[26 +: 1]),

    .AXI_26_ARADDR(m_axi_hbm_int_araddr[26*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_26_ARBURST(m_axi_hbm_int_arburst[26*2 +: 2]),
    .AXI_26_ARID(m_axi_hbm_int_arid[26*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_26_ARLEN(m_axi_hbm_int_arlen[26*8 +: 4]),
    .AXI_26_ARSIZE(m_axi_hbm_int_arsize[26*3 +: 3]),
    .AXI_26_ARVALID(m_axi_hbm_int_arvalid[26 +: 1]),
    .AXI_26_ARREADY(m_axi_hbm_int_arready[26 +: 1]),
    .AXI_26_RDATA_PARITY(),
    .AXI_26_RDATA(m_axi_hbm_int_rdata[26*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_26_RID(m_axi_hbm_int_rid[26*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_26_RLAST(m_axi_hbm_int_rlast[26 +: 1]),
    .AXI_26_RRESP(m_axi_hbm_int_rresp[26*2 +: 2]),
    .AXI_26_RVALID(m_axi_hbm_int_rvalid[26 +: 1]),
    .AXI_26_RREADY(m_axi_hbm_int_rready[26 +: 1]),
    .AXI_26_AWADDR(m_axi_hbm_int_awaddr[26*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_26_AWBURST(m_axi_hbm_int_awburst[26*2 +: 2]),
    .AXI_26_AWID(m_axi_hbm_int_awid[26*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_26_AWLEN(m_axi_hbm_int_awlen[26*8 +: 4]),
    .AXI_26_AWSIZE(m_axi_hbm_int_awsize[26*3 +: 3]),
    .AXI_26_AWVALID(m_axi_hbm_int_awvalid[26 +: 1]),
    .AXI_26_AWREADY(m_axi_hbm_int_awready[26 +: 1]),
    .AXI_26_WDATA(m_axi_hbm_int_wdata[26*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_26_WLAST(m_axi_hbm_int_wlast[26 +: 1]),
    .AXI_26_WSTRB(m_axi_hbm_int_wstrb[26*AXI_HBM_STRB_WIDTH +: AXI_HBM_STRB_WIDTH]),
    .AXI_26_WDATA_PARITY(32'd0),
    .AXI_26_WVALID(m_axi_hbm_int_wvalid[26 +: 1]),
    .AXI_26_WREADY(m_axi_hbm_int_wready[26 +: 1]),
    .AXI_26_BID(m_axi_hbm_int_bid[26*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_26_BRESP(m_axi_hbm_int_bresp[26*2 +: 2]),
    .AXI_26_BVALID(m_axi_hbm_int_bvalid[26 +: 1]),
    .AXI_26_BREADY(m_axi_hbm_int_bready[26 +: 1]),

    .AXI_27_ACLK(hbm_clk_int[27 +: 1]),
    .AXI_27_ARESET_N(!hbm_rst_int[27 +: 1]),

    .AXI_27_ARADDR(m_axi_hbm_int_araddr[27*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_27_ARBURST(m_axi_hbm_int_arburst[27*2 +: 2]),
    .AXI_27_ARID(m_axi_hbm_int_arid[27*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_27_ARLEN(m_axi_hbm_int_arlen[27*8 +: 4]),
    .AXI_27_ARSIZE(m_axi_hbm_int_arsize[27*3 +: 3]),
    .AXI_27_ARVALID(m_axi_hbm_int_arvalid[27 +: 1]),
    .AXI_27_ARREADY(m_axi_hbm_int_arready[27 +: 1]),
    .AXI_27_RDATA_PARITY(),
    .AXI_27_RDATA(m_axi_hbm_int_rdata[27*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_27_RID(m_axi_hbm_int_rid[27*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_27_RLAST(m_axi_hbm_int_rlast[27 +: 1]),
    .AXI_27_RRESP(m_axi_hbm_int_rresp[27*2 +: 2]),
    .AXI_27_RVALID(m_axi_hbm_int_rvalid[27 +: 1]),
    .AXI_27_RREADY(m_axi_hbm_int_rready[27 +: 1]),
    .AXI_27_AWADDR(m_axi_hbm_int_awaddr[27*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_27_AWBURST(m_axi_hbm_int_awburst[27*2 +: 2]),
    .AXI_27_AWID(m_axi_hbm_int_awid[27*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_27_AWLEN(m_axi_hbm_int_awlen[27*8 +: 4]),
    .AXI_27_AWSIZE(m_axi_hbm_int_awsize[27*3 +: 3]),
    .AXI_27_AWVALID(m_axi_hbm_int_awvalid[27 +: 1]),
    .AXI_27_AWREADY(m_axi_hbm_int_awready[27 +: 1]),
    .AXI_27_WDATA(m_axi_hbm_int_wdata[27*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_27_WLAST(m_axi_hbm_int_wlast[27 +: 1]),
    .AXI_27_WSTRB(m_axi_hbm_int_wstrb[27*AXI_HBM_STRB_WIDTH +: AXI_HBM_STRB_WIDTH]),
    .AXI_27_WDATA_PARITY(32'd0),
    .AXI_27_WVALID(m_axi_hbm_int_wvalid[27 +: 1]),
    .AXI_27_WREADY(m_axi_hbm_int_wready[27 +: 1]),
    .AXI_27_BID(m_axi_hbm_int_bid[27*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_27_BRESP(m_axi_hbm_int_bresp[27*2 +: 2]),
    .AXI_27_BVALID(m_axi_hbm_int_bvalid[27 +: 1]),
    .AXI_27_BREADY(m_axi_hbm_int_bready[27 +: 1]),

    .AXI_28_ACLK(hbm_clk_int[28 +: 1]),
    .AXI_28_ARESET_N(!hbm_rst_int[28 +: 1]),

    .AXI_28_ARADDR(m_axi_hbm_int_araddr[28*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_28_ARBURST(m_axi_hbm_int_arburst[28*2 +: 2]),
    .AXI_28_ARID(m_axi_hbm_int_arid[28*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_28_ARLEN(m_axi_hbm_int_arlen[28*8 +: 4]),
    .AXI_28_ARSIZE(m_axi_hbm_int_arsize[28*3 +: 3]),
    .AXI_28_ARVALID(m_axi_hbm_int_arvalid[28 +: 1]),
    .AXI_28_ARREADY(m_axi_hbm_int_arready[28 +: 1]),
    .AXI_28_RDATA_PARITY(),
    .AXI_28_RDATA(m_axi_hbm_int_rdata[28*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_28_RID(m_axi_hbm_int_rid[28*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_28_RLAST(m_axi_hbm_int_rlast[28 +: 1]),
    .AXI_28_RRESP(m_axi_hbm_int_rresp[28*2 +: 2]),
    .AXI_28_RVALID(m_axi_hbm_int_rvalid[28 +: 1]),
    .AXI_28_RREADY(m_axi_hbm_int_rready[28 +: 1]),
    .AXI_28_AWADDR(m_axi_hbm_int_awaddr[28*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_28_AWBURST(m_axi_hbm_int_awburst[28*2 +: 2]),
    .AXI_28_AWID(m_axi_hbm_int_awid[28*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_28_AWLEN(m_axi_hbm_int_awlen[28*8 +: 4]),
    .AXI_28_AWSIZE(m_axi_hbm_int_awsize[28*3 +: 3]),
    .AXI_28_AWVALID(m_axi_hbm_int_awvalid[28 +: 1]),
    .AXI_28_AWREADY(m_axi_hbm_int_awready[28 +: 1]),
    .AXI_28_WDATA(m_axi_hbm_int_wdata[28*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_28_WLAST(m_axi_hbm_int_wlast[28 +: 1]),
    .AXI_28_WSTRB(m_axi_hbm_int_wstrb[28*AXI_HBM_STRB_WIDTH +: AXI_HBM_STRB_WIDTH]),
    .AXI_28_WDATA_PARITY(32'd0),
    .AXI_28_WVALID(m_axi_hbm_int_wvalid[28 +: 1]),
    .AXI_28_WREADY(m_axi_hbm_int_wready[28 +: 1]),
    .AXI_28_BID(m_axi_hbm_int_bid[28*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_28_BRESP(m_axi_hbm_int_bresp[28*2 +: 2]),
    .AXI_28_BVALID(m_axi_hbm_int_bvalid[28 +: 1]),
    .AXI_28_BREADY(m_axi_hbm_int_bready[28 +: 1]),

    .AXI_29_ACLK(hbm_clk_int[29 +: 1]),
    .AXI_29_ARESET_N(!hbm_rst_int[29 +: 1]),

    .AXI_29_ARADDR(m_axi_hbm_int_araddr[29*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_29_ARBURST(m_axi_hbm_int_arburst[29*2 +: 2]),
    .AXI_29_ARID(m_axi_hbm_int_arid[29*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_29_ARLEN(m_axi_hbm_int_arlen[29*8 +: 4]),
    .AXI_29_ARSIZE(m_axi_hbm_int_arsize[29*3 +: 3]),
    .AXI_29_ARVALID(m_axi_hbm_int_arvalid[29 +: 1]),
    .AXI_29_ARREADY(m_axi_hbm_int_arready[29 +: 1]),
    .AXI_29_RDATA_PARITY(),
    .AXI_29_RDATA(m_axi_hbm_int_rdata[29*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_29_RID(m_axi_hbm_int_rid[29*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_29_RLAST(m_axi_hbm_int_rlast[29 +: 1]),
    .AXI_29_RRESP(m_axi_hbm_int_rresp[29*2 +: 2]),
    .AXI_29_RVALID(m_axi_hbm_int_rvalid[29 +: 1]),
    .AXI_29_RREADY(m_axi_hbm_int_rready[29 +: 1]),
    .AXI_29_AWADDR(m_axi_hbm_int_awaddr[29*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_29_AWBURST(m_axi_hbm_int_awburst[29*2 +: 2]),
    .AXI_29_AWID(m_axi_hbm_int_awid[29*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_29_AWLEN(m_axi_hbm_int_awlen[29*8 +: 4]),
    .AXI_29_AWSIZE(m_axi_hbm_int_awsize[29*3 +: 3]),
    .AXI_29_AWVALID(m_axi_hbm_int_awvalid[29 +: 1]),
    .AXI_29_AWREADY(m_axi_hbm_int_awready[29 +: 1]),
    .AXI_29_WDATA(m_axi_hbm_int_wdata[29*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_29_WLAST(m_axi_hbm_int_wlast[29 +: 1]),
    .AXI_29_WSTRB(m_axi_hbm_int_wstrb[29*AXI_HBM_STRB_WIDTH +: AXI_HBM_STRB_WIDTH]),
    .AXI_29_WDATA_PARITY(32'd0),
    .AXI_29_WVALID(m_axi_hbm_int_wvalid[29 +: 1]),
    .AXI_29_WREADY(m_axi_hbm_int_wready[29 +: 1]),
    .AXI_29_BID(m_axi_hbm_int_bid[29*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_29_BRESP(m_axi_hbm_int_bresp[29*2 +: 2]),
    .AXI_29_BVALID(m_axi_hbm_int_bvalid[29 +: 1]),
    .AXI_29_BREADY(m_axi_hbm_int_bready[29 +: 1]),

    .AXI_30_ACLK(hbm_clk_int[30 +: 1]),
    .AXI_30_ARESET_N(!hbm_rst_int[30 +: 1]),

    .AXI_30_ARADDR(m_axi_hbm_int_araddr[30*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_30_ARBURST(m_axi_hbm_int_arburst[30*2 +: 2]),
    .AXI_30_ARID(m_axi_hbm_int_arid[30*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_30_ARLEN(m_axi_hbm_int_arlen[30*8 +: 4]),
    .AXI_30_ARSIZE(m_axi_hbm_int_arsize[30*3 +: 3]),
    .AXI_30_ARVALID(m_axi_hbm_int_arvalid[30 +: 1]),
    .AXI_30_ARREADY(m_axi_hbm_int_arready[30 +: 1]),
    .AXI_30_RDATA_PARITY(),
    .AXI_30_RDATA(m_axi_hbm_int_rdata[30*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_30_RID(m_axi_hbm_int_rid[30*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_30_RLAST(m_axi_hbm_int_rlast[30 +: 1]),
    .AXI_30_RRESP(m_axi_hbm_int_rresp[30*2 +: 2]),
    .AXI_30_RVALID(m_axi_hbm_int_rvalid[30 +: 1]),
    .AXI_30_RREADY(m_axi_hbm_int_rready[30 +: 1]),
    .AXI_30_AWADDR(m_axi_hbm_int_awaddr[30*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_30_AWBURST(m_axi_hbm_int_awburst[30*2 +: 2]),
    .AXI_30_AWID(m_axi_hbm_int_awid[30*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_30_AWLEN(m_axi_hbm_int_awlen[30*8 +: 4]),
    .AXI_30_AWSIZE(m_axi_hbm_int_awsize[30*3 +: 3]),
    .AXI_30_AWVALID(m_axi_hbm_int_awvalid[30 +: 1]),
    .AXI_30_AWREADY(m_axi_hbm_int_awready[30 +: 1]),
    .AXI_30_WDATA(m_axi_hbm_int_wdata[30*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_30_WLAST(m_axi_hbm_int_wlast[30 +: 1]),
    .AXI_30_WSTRB(m_axi_hbm_int_wstrb[30*AXI_HBM_STRB_WIDTH +: AXI_HBM_STRB_WIDTH]),
    .AXI_30_WDATA_PARITY(32'd0),
    .AXI_30_WVALID(m_axi_hbm_int_wvalid[30 +: 1]),
    .AXI_30_WREADY(m_axi_hbm_int_wready[30 +: 1]),
    .AXI_30_BID(m_axi_hbm_int_bid[30*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_30_BRESP(m_axi_hbm_int_bresp[30*2 +: 2]),
    .AXI_30_BVALID(m_axi_hbm_int_bvalid[30 +: 1]),
    .AXI_30_BREADY(m_axi_hbm_int_bready[30 +: 1]),

    .AXI_31_ACLK(hbm_clk_int[31 +: 1]),
    .AXI_31_ARESET_N(!hbm_rst_int[31 +: 1]),

    .AXI_31_ARADDR(m_axi_hbm_int_araddr[31*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_31_ARBURST(m_axi_hbm_int_arburst[31*2 +: 2]),
    .AXI_31_ARID(m_axi_hbm_int_arid[31*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_31_ARLEN(m_axi_hbm_int_arlen[31*8 +: 4]),
    .AXI_31_ARSIZE(m_axi_hbm_int_arsize[31*3 +: 3]),
    .AXI_31_ARVALID(m_axi_hbm_int_arvalid[31 +: 1]),
    .AXI_31_ARREADY(m_axi_hbm_int_arready[31 +: 1]),
    .AXI_31_RDATA_PARITY(),
    .AXI_31_RDATA(m_axi_hbm_int_rdata[31*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_31_RID(m_axi_hbm_int_rid[31*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_31_RLAST(m_axi_hbm_int_rlast[31 +: 1]),
    .AXI_31_RRESP(m_axi_hbm_int_rresp[31*2 +: 2]),
    .AXI_31_RVALID(m_axi_hbm_int_rvalid[31 +: 1]),
    .AXI_31_RREADY(m_axi_hbm_int_rready[31 +: 1]),
    .AXI_31_AWADDR(m_axi_hbm_int_awaddr[31*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH]),
    .AXI_31_AWBURST(m_axi_hbm_int_awburst[31*2 +: 2]),
    .AXI_31_AWID(m_axi_hbm_int_awid[31*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_31_AWLEN(m_axi_hbm_int_awlen[31*8 +: 4]),
    .AXI_31_AWSIZE(m_axi_hbm_int_awsize[31*3 +: 3]),
    .AXI_31_AWVALID(m_axi_hbm_int_awvalid[31 +: 1]),
    .AXI_31_AWREADY(m_axi_hbm_int_awready[31 +: 1]),
    .AXI_31_WDATA(m_axi_hbm_int_wdata[31*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH]),
    .AXI_31_WLAST(m_axi_hbm_int_wlast[31 +: 1]),
    .AXI_31_WSTRB(m_axi_hbm_int_wstrb[31*AXI_HBM_STRB_WIDTH +: AXI_HBM_STRB_WIDTH]),
    .AXI_31_WDATA_PARITY(32'd0),
    .AXI_31_WVALID(m_axi_hbm_int_wvalid[31 +: 1]),
    .AXI_31_WREADY(m_axi_hbm_int_wready[31 +: 1]),
    .AXI_31_BID(m_axi_hbm_int_bid[31*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH]),
    .AXI_31_BRESP(m_axi_hbm_int_bresp[31*2 +: 2]),
    .AXI_31_BVALID(m_axi_hbm_int_bvalid[31 +: 1]),
    .AXI_31_BREADY(m_axi_hbm_int_bready[31 +: 1]),

    .DRAM_0_STAT_CATTRIP(hbm_cattrip_1),
    .DRAM_0_STAT_TEMP(hbm_temp_1),
    .DRAM_1_STAT_CATTRIP(hbm_cattrip_2),
    .DRAM_1_STAT_TEMP(hbm_temp_2)
);

for (n = 0; n < HBM_CH_INT; n = n + 1) begin

    localparam c = n / HBM_CH_STRIDE;

    if (c*HBM_CH_STRIDE == n) begin

        assign hbm_clk[c] = hbm_clk_int[n];
        assign hbm_rst[c] = hbm_rst_int[n];

        assign m_axi_hbm_int_awid[n*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH] = s_axi_hbm_awid[c*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH];
        assign m_axi_hbm_int_awaddr[n*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH] = s_axi_hbm_awaddr[c*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH];
        assign m_axi_hbm_int_awlen[n*8 +: 8] = s_axi_hbm_awlen[c*8 +: 8];
        assign m_axi_hbm_int_awsize[n*3 +: 3] = s_axi_hbm_awsize[c*3 +: 3];
        assign m_axi_hbm_int_awburst[n*2 +: 2] = s_axi_hbm_awburst[c*2 +: 2];
        assign m_axi_hbm_int_awlock[n*1 +: 1] = s_axi_hbm_awlock[c*1 +: 1];
        assign m_axi_hbm_int_awcache[n*4 +: 4] = s_axi_hbm_awcache[c*4 +: 4];
        assign m_axi_hbm_int_awprot[n*3 +: 3] = s_axi_hbm_awprot[c*3 +: 3];
        assign m_axi_hbm_int_awqos[n*4 +: 4] = s_axi_hbm_awqos[c*4 +: 4];
        assign m_axi_hbm_int_awvalid[n*1 +: 1] = s_axi_hbm_awvalid[c*1 +: 1];
        assign s_axi_hbm_awready[c*1 +: 1] = m_axi_hbm_int_awready[n*1 +: 1];
        assign m_axi_hbm_int_wdata[n*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH] = s_axi_hbm_wdata[c*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH];
        assign m_axi_hbm_int_wstrb[n*AXI_HBM_STRB_WIDTH +: AXI_HBM_STRB_WIDTH] = s_axi_hbm_wstrb[c*AXI_HBM_STRB_WIDTH +: AXI_HBM_STRB_WIDTH];
        assign m_axi_hbm_int_wlast[n*1 +: 1] = s_axi_hbm_wlast[c*1 +: 1];
        assign m_axi_hbm_int_wvalid[n*1 +: 1] = s_axi_hbm_wvalid[c*1 +: 1];
        assign s_axi_hbm_wready[c*1 +: 1] = m_axi_hbm_int_wready[n*1 +: 1];
        assign s_axi_hbm_bid[c*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH] = m_axi_hbm_int_bid[n*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH];
        assign s_axi_hbm_bresp[c*2 +: 2] = m_axi_hbm_int_bresp[n*2 +: 2];
        assign s_axi_hbm_bvalid[c*1 +: 1] = m_axi_hbm_int_bvalid[n*1 +: 1];
        assign m_axi_hbm_int_bready[n*1 +: 1] = s_axi_hbm_bready[c*1 +: 1];
        assign m_axi_hbm_int_arid[n*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH] = s_axi_hbm_arid[c*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH];
        assign m_axi_hbm_int_araddr[n*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH] = s_axi_hbm_araddr[c*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH];
        assign m_axi_hbm_int_arlen[n*8 +: 8] = s_axi_hbm_arlen[c*8 +: 8];
        assign m_axi_hbm_int_arsize[n*3 +: 3] = s_axi_hbm_arsize[c*3 +: 3];
        assign m_axi_hbm_int_arburst[n*2 +: 2] = s_axi_hbm_arburst[c*2 +: 2];
        assign m_axi_hbm_int_arlock[n*1 +: 1] = s_axi_hbm_arlock[c*1 +: 1];
        assign m_axi_hbm_int_arcache[n*4 +: 4] = s_axi_hbm_arcache[c*4 +: 4];
        assign m_axi_hbm_int_arprot[n*3 +: 3] = s_axi_hbm_arprot[c*3 +: 3];
        assign m_axi_hbm_int_arqos[n*4 +: 4] = s_axi_hbm_arqos[c*4 +: 4];
        assign m_axi_hbm_int_arvalid[n*1 +: 1] = s_axi_hbm_arvalid[c*1 +: 1];
        assign s_axi_hbm_arready[c*1 +: 1] = m_axi_hbm_int_arready[n*1 +: 1];
        assign s_axi_hbm_rid[c*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH] = m_axi_hbm_int_rid[n*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH];
        assign s_axi_hbm_rdata[c*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH] = m_axi_hbm_int_rdata[n*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH];
        assign s_axi_hbm_rresp[c*2 +: 2] = m_axi_hbm_int_rresp[n*2 +: 2];
        assign s_axi_hbm_rlast[c*1 +: 1] = m_axi_hbm_int_rlast[n*1 +: 1];
        assign s_axi_hbm_rvalid[c*1 +: 1] = m_axi_hbm_int_rvalid[n*1 +: 1];
        assign m_axi_hbm_int_rready[n*1 +: 1] = s_axi_hbm_rready[c*1 +: 1];

        assign hbm_status[c] = !hbm_rst_int[n];

    end else begin

        assign m_axi_hbm_int_awid[n*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH] = 0;
        assign m_axi_hbm_int_awaddr[n*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH] = 0;
        assign m_axi_hbm_int_awlen[n*8 +: 8] = 8'd0;
        assign m_axi_hbm_int_awsize[n*3 +: 3] = 3'd0;
        assign m_axi_hbm_int_awburst[n*2 +: 2] = 2'd0;
        assign m_axi_hbm_int_awlock[n*1 +: 1] = 1'b0;
        assign m_axi_hbm_int_awcache[n*4 +: 4] = 4'd0;
        assign m_axi_hbm_int_awprot[n*3 +: 3] = 3'd0;
        assign m_axi_hbm_int_awqos[n*4 +: 4] = 4'd0;
        assign m_axi_hbm_int_awvalid[n*1 +: 1] = 1'b0;
        assign m_axi_hbm_int_wdata[n*AXI_HBM_DATA_WIDTH +: AXI_HBM_DATA_WIDTH] = 0;
        assign m_axi_hbm_int_wstrb[n*AXI_HBM_STRB_WIDTH +: AXI_HBM_STRB_WIDTH] = 0;
        assign m_axi_hbm_int_wlast[n*1 +: 1] = 1'b0;
        assign m_axi_hbm_int_wvalid[n*1 +: 1] = 1'b0;
        assign m_axi_hbm_int_bready[n*1 +: 1] = 1'b1;
        assign m_axi_hbm_int_arid[n*AXI_HBM_ID_WIDTH +: AXI_HBM_ID_WIDTH] = 0;
        assign m_axi_hbm_int_araddr[n*AXI_HBM_ADDR_WIDTH +: AXI_HBM_ADDR_WIDTH] = 0;
        assign m_axi_hbm_int_arlen[n*8 +: 8] = 8'd0;
        assign m_axi_hbm_int_arsize[n*3 +: 3] = 3'd0;
        assign m_axi_hbm_int_arburst[n*2 +: 2] = 2'd0;
        assign m_axi_hbm_int_arlock[n*1 +: 1] = 1'b0;
        assign m_axi_hbm_int_arcache[n*4 +: 4] = 4'd0;
        assign m_axi_hbm_int_arprot[n*3 +: 3] = 3'd0;
        assign m_axi_hbm_int_arqos[n*4 +: 4] = 4'd0;
        assign m_axi_hbm_int_arvalid[n*1 +: 1] = 1'b0;
        assign m_axi_hbm_int_rready[n*1 +: 1] = 1'b1;

    end

end

endgenerate

endmodule

`resetall
